module s27(input clk,input in[9:0], output out);
reg[2:0] state;
