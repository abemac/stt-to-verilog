module s820(input clk,input[9:0] in, output [7:0] out);
	reg[4:0] state;
	always @(posedge clk) begin
		out<=0;
		case (state)
			0: begin
				if(in == 0) begin
					state<=1;
					out<=0;
				end
			end
			1: begin
				if(in == 0) begin
					state<=1;
					out<=1;
				end
				if(in == 1) begin
					state<=1;
					out<=2;
				end
				if(in == 2) begin
					state<=17;
					out<=3;
				end
				if(in == 3) begin
					state<=1;
					out<=4;
				end
				if(in == 4) begin
					state<=17;
					out<=5;
				end
				if(in == 5) begin
					state<=1;
					out<=6;
				end
				if(in == 6) begin
					state<=17;
					out<=7;
				end
				if(in == 7) begin
					state<=17;
					out<=8;
				end
				if(in == 8) begin
					state<=17;
					out<=9;
				end
				if(in == 9) begin
					state<=17;
					out<=10;
				end
				if(in == 10) begin
					state<=17;
					out<=11;
				end
				if(in == 11) begin
					state<=17;
					out<=12;
				end
				if(in == 12) begin
					state<=17;
					out<=13;
				end
				if(in == 13) begin
					state<=17;
					out<=14;
				end
				if(in == 14) begin
					state<=17;
					out<=15;
				end
				if(in == 15) begin
					state<=17;
					out<=16;
				end
				if(in == 16) begin
					state<=17;
					out<=17;
				end
				if(in == 17) begin
					state<=17;
					out<=18;
				end
				if(in == 18) begin
					state<=17;
					out<=19;
				end
				if(in == 19) begin
					state<=17;
					out<=20;
				end
				if(in == 20) begin
					state<=17;
					out<=21;
				end
				if(in == 21) begin
					state<=17;
					out<=22;
				end
				if(in == 22) begin
					state<=17;
					out<=23;
				end
				if(in == 23) begin
					state<=17;
					out<=24;
				end
				if(in == 24) begin
					state<=17;
					out<=25;
				end
				if(in == 25) begin
					state<=17;
					out<=26;
				end
				if(in == 26) begin
					state<=17;
					out<=27;
				end
				if(in == 27) begin
					state<=17;
					out<=28;
				end
				if(in == 28) begin
					state<=17;
					out<=29;
				end
				if(in == 29) begin
					state<=17;
					out<=30;
				end
				if(in == 30) begin
					state<=17;
					out<=31;
				end
				if(in == 31) begin
					state<=17;
					out<=32;
				end
				if(in == 32) begin
					state<=17;
					out<=33;
				end
				if(in == 33) begin
					state<=17;
					out<=34;
				end
				if(in == 34) begin
					state<=17;
					out<=35;
				end
				if(in == 35) begin
					state<=17;
					out<=36;
				end
				if(in == 36) begin
					state<=17;
					out<=37;
				end
				if(in == 37) begin
					state<=17;
					out<=38;
				end
				if(in == 38) begin
					state<=17;
					out<=39;
				end
				if(in == 39) begin
					state<=17;
					out<=40;
				end
				if(in == 40) begin
					state<=17;
					out<=41;
				end
				if(in == 41) begin
					state<=17;
					out<=42;
				end
				if(in == 42) begin
					state<=17;
					out<=43;
				end
				if(in == 43) begin
					state<=17;
					out<=44;
				end
				if(in == 44) begin
					state<=17;
					out<=45;
				end
				if(in == 45) begin
					state<=17;
					out<=46;
				end
				if(in == 46) begin
					state<=17;
					out<=47;
				end
				if(in == 47) begin
					state<=17;
					out<=48;
				end
				if(in == 48) begin
					state<=17;
					out<=49;
				end
				if(in == 49) begin
					state<=17;
					out<=50;
				end
				if(in == 50) begin
					state<=17;
					out<=51;
				end
				if(in == 51) begin
					state<=17;
					out<=52;
				end
				if(in == 52) begin
					state<=17;
					out<=53;
				end
				if(in == 53) begin
					state<=1;
					out<=54;
				end
				if(in == 54) begin
					state<=17;
					out<=55;
				end
				if(in == 55) begin
					state<=1;
					out<=56;
				end
				if(in == 56) begin
					state<=17;
					out<=57;
				end
				if(in == 57) begin
					state<=1;
					out<=58;
				end
				if(in == 58) begin
					state<=17;
					out<=59;
				end
				if(in == 59) begin
					state<=17;
					out<=60;
				end
				if(in == 60) begin
					state<=17;
					out<=61;
				end
				if(in == 61) begin
					state<=17;
					out<=62;
				end
				if(in == 62) begin
					state<=17;
					out<=63;
				end
				if(in == 63) begin
					state<=17;
					out<=64;
				end
				if(in == 64) begin
					state<=17;
					out<=65;
				end
				if(in == 65) begin
					state<=17;
					out<=66;
				end
				if(in == 66) begin
					state<=17;
					out<=67;
				end
				if(in == 67) begin
					state<=17;
					out<=68;
				end
				if(in == 68) begin
					state<=17;
					out<=69;
				end
				if(in == 69) begin
					state<=17;
					out<=70;
				end
				if(in == 70) begin
					state<=17;
					out<=71;
				end
				if(in == 71) begin
					state<=17;
					out<=72;
				end
				if(in == 72) begin
					state<=17;
					out<=73;
				end
				if(in == 73) begin
					state<=17;
					out<=74;
				end
				if(in == 74) begin
					state<=17;
					out<=75;
				end
				if(in == 75) begin
					state<=17;
					out<=76;
				end
				if(in == 76) begin
					state<=17;
					out<=77;
				end
				if(in == 77) begin
					state<=17;
					out<=78;
				end
				if(in == 78) begin
					state<=17;
					out<=79;
				end
				if(in == 79) begin
					state<=17;
					out<=80;
				end
				if(in == 80) begin
					state<=17;
					out<=81;
				end
				if(in == 81) begin
					state<=17;
					out<=82;
				end
				if(in == 82) begin
					state<=17;
					out<=83;
				end
				if(in == 83) begin
					state<=17;
					out<=84;
				end
				if(in == 84) begin
					state<=17;
					out<=85;
				end
				if(in == 85) begin
					state<=17;
					out<=86;
				end
				if(in == 86) begin
					state<=17;
					out<=87;
				end
				if(in == 87) begin
					state<=17;
					out<=88;
				end
				if(in == 88) begin
					state<=17;
					out<=89;
				end
				if(in == 89) begin
					state<=17;
					out<=90;
				end
				if(in == 90) begin
					state<=17;
					out<=91;
				end
				if(in == 91) begin
					state<=17;
					out<=92;
				end
				if(in == 92) begin
					state<=17;
					out<=93;
				end
				if(in == 93) begin
					state<=17;
					out<=94;
				end
				if(in == 94) begin
					state<=17;
					out<=95;
				end
				if(in == 95) begin
					state<=17;
					out<=96;
				end
				if(in == 96) begin
					state<=17;
					out<=97;
				end
				if(in == 97) begin
					state<=17;
					out<=98;
				end
				if(in == 98) begin
					state<=17;
					out<=99;
				end
				if(in == 99) begin
					state<=17;
					out<=100;
				end
				if(in == 100) begin
					state<=17;
					out<=101;
				end
				if(in == 101) begin
					state<=17;
					out<=102;
				end
				if(in == 102) begin
					state<=17;
					out<=103;
				end
				if(in == 103) begin
					state<=17;
					out<=104;
				end
				if(in == 104) begin
					state<=17;
					out<=105;
				end
				if(in == 105) begin
					state<=1;
					out<=106;
				end
				if(in == 106) begin
					state<=17;
					out<=107;
				end
				if(in == 107) begin
					state<=1;
					out<=108;
				end
				if(in == 108) begin
					state<=17;
					out<=109;
				end
				if(in == 109) begin
					state<=1;
					out<=110;
				end
				if(in == 110) begin
					state<=17;
					out<=111;
				end
				if(in == 111) begin
					state<=1;
					out<=112;
				end
				if(in == 112) begin
					state<=17;
					out<=113;
				end
				if(in == 113) begin
					state<=1;
					out<=114;
				end
				if(in == 114) begin
					state<=17;
					out<=115;
				end
				if(in == 115) begin
					state<=1;
					out<=116;
				end
				if(in == 116) begin
					state<=17;
					out<=117;
				end
				if(in == 117) begin
					state<=1;
					out<=118;
				end
				if(in == 118) begin
					state<=17;
					out<=119;
				end
				if(in == 119) begin
					state<=1;
					out<=120;
				end
				if(in == 120) begin
					state<=17;
					out<=121;
				end
				if(in == 121) begin
					state<=1;
					out<=122;
				end
				if(in == 122) begin
					state<=17;
					out<=123;
				end
				if(in == 123) begin
					state<=17;
					out<=124;
				end
				if(in == 124) begin
					state<=17;
					out<=125;
				end
				if(in == 125) begin
					state<=17;
					out<=126;
				end
				if(in == 126) begin
					state<=17;
					out<=127;
				end
				if(in == 127) begin
					state<=17;
					out<=128;
				end
				if(in == 128) begin
					state<=17;
					out<=129;
				end
				if(in == 129) begin
					state<=17;
					out<=130;
				end
				if(in == 130) begin
					state<=17;
					out<=131;
				end
				if(in == 131) begin
					state<=17;
					out<=132;
				end
				if(in == 132) begin
					state<=17;
					out<=133;
				end
				if(in == 133) begin
					state<=17;
					out<=134;
				end
				if(in == 134) begin
					state<=17;
					out<=135;
				end
				if(in == 135) begin
					state<=17;
					out<=136;
				end
				if(in == 136) begin
					state<=17;
					out<=137;
				end
				if(in == 137) begin
					state<=17;
					out<=138;
				end
				if(in == 138) begin
					state<=17;
					out<=139;
				end
				if(in == 139) begin
					state<=17;
					out<=140;
				end
				if(in == 140) begin
					state<=17;
					out<=141;
				end
				if(in == 141) begin
					state<=17;
					out<=142;
				end
				if(in == 142) begin
					state<=17;
					out<=143;
				end
				if(in == 143) begin
					state<=17;
					out<=144;
				end
				if(in == 144) begin
					state<=17;
					out<=145;
				end
				if(in == 145) begin
					state<=17;
					out<=146;
				end
				if(in == 146) begin
					state<=17;
					out<=147;
				end
				if(in == 147) begin
					state<=17;
					out<=148;
				end
				if(in == 148) begin
					state<=17;
					out<=149;
				end
				if(in == 149) begin
					state<=17;
					out<=150;
				end
				if(in == 150) begin
					state<=17;
					out<=151;
				end
				if(in == 151) begin
					state<=17;
					out<=152;
				end
				if(in == 152) begin
					state<=17;
					out<=153;
				end
				if(in == 153) begin
					state<=17;
					out<=154;
				end
				if(in == 154) begin
					state<=17;
					out<=155;
				end
				if(in == 155) begin
					state<=17;
					out<=156;
				end
				if(in == 156) begin
					state<=17;
					out<=157;
				end
				if(in == 157) begin
					state<=17;
					out<=158;
				end
				if(in == 158) begin
					state<=17;
					out<=159;
				end
				if(in == 159) begin
					state<=17;
					out<=160;
				end
				if(in == 160) begin
					state<=17;
					out<=161;
				end
				if(in == 161) begin
					state<=17;
					out<=162;
				end
				if(in == 162) begin
					state<=17;
					out<=163;
				end
				if(in == 163) begin
					state<=17;
					out<=164;
				end
				if(in == 164) begin
					state<=17;
					out<=165;
				end
				if(in == 165) begin
					state<=17;
					out<=166;
				end
				if(in == 166) begin
					state<=17;
					out<=167;
				end
				if(in == 167) begin
					state<=17;
					out<=168;
				end
				if(in == 168) begin
					state<=17;
					out<=169;
				end
				if(in == 169) begin
					state<=1;
					out<=170;
				end
				if(in == 170) begin
					state<=17;
					out<=171;
				end
				if(in == 171) begin
					state<=1;
					out<=172;
				end
				if(in == 172) begin
					state<=17;
					out<=173;
				end
				if(in == 173) begin
					state<=1;
					out<=174;
				end
				if(in == 174) begin
					state<=17;
					out<=175;
				end
				if(in == 175) begin
					state<=17;
					out<=176;
				end
				if(in == 176) begin
					state<=17;
					out<=177;
				end
				if(in == 177) begin
					state<=17;
					out<=178;
				end
				if(in == 178) begin
					state<=17;
					out<=179;
				end
				if(in == 179) begin
					state<=17;
					out<=180;
				end
				if(in == 180) begin
					state<=17;
					out<=181;
				end
				if(in == 181) begin
					state<=17;
					out<=182;
				end
				if(in == 182) begin
					state<=17;
					out<=183;
				end
				if(in == 183) begin
					state<=17;
					out<=184;
				end
				if(in == 184) begin
					state<=17;
					out<=185;
				end
				if(in == 185) begin
					state<=17;
					out<=186;
				end
				if(in == 186) begin
					state<=17;
					out<=187;
				end
				if(in == 187) begin
					state<=17;
					out<=188;
				end
				if(in == 188) begin
					state<=17;
					out<=189;
				end
				if(in == 189) begin
					state<=17;
					out<=190;
				end
				if(in == 190) begin
					state<=17;
					out<=191;
				end
				if(in == 191) begin
					state<=17;
					out<=192;
				end
				if(in == 192) begin
					state<=17;
					out<=193;
				end
				if(in == 193) begin
					state<=17;
					out<=194;
				end
				if(in == 194) begin
					state<=17;
					out<=195;
				end
				if(in == 195) begin
					state<=17;
					out<=196;
				end
				if(in == 196) begin
					state<=17;
					out<=197;
				end
				if(in == 197) begin
					state<=17;
					out<=198;
				end
				if(in == 198) begin
					state<=17;
					out<=199;
				end
				if(in == 199) begin
					state<=17;
					out<=200;
				end
				if(in == 200) begin
					state<=17;
					out<=201;
				end
				if(in == 201) begin
					state<=17;
					out<=202;
				end
				if(in == 202) begin
					state<=17;
					out<=203;
				end
				if(in == 203) begin
					state<=17;
					out<=204;
				end
				if(in == 204) begin
					state<=17;
					out<=205;
				end
				if(in == 205) begin
					state<=17;
					out<=206;
				end
				if(in == 206) begin
					state<=17;
					out<=207;
				end
				if(in == 207) begin
					state<=17;
					out<=208;
				end
				if(in == 208) begin
					state<=17;
					out<=209;
				end
				if(in == 209) begin
					state<=17;
					out<=210;
				end
				if(in == 210) begin
					state<=17;
					out<=211;
				end
				if(in == 211) begin
					state<=17;
					out<=212;
				end
				if(in == 212) begin
					state<=17;
					out<=213;
				end
				if(in == 213) begin
					state<=17;
					out<=214;
				end
				if(in == 214) begin
					state<=17;
					out<=215;
				end
				if(in == 215) begin
					state<=17;
					out<=216;
				end
				if(in == 216) begin
					state<=17;
					out<=217;
				end
				if(in == 217) begin
					state<=17;
					out<=218;
				end
				if(in == 218) begin
					state<=17;
					out<=219;
				end
				if(in == 219) begin
					state<=17;
					out<=220;
				end
				if(in == 220) begin
					state<=17;
					out<=221;
				end
				if(in == 221) begin
					state<=1;
					out<=222;
				end
				if(in == 222) begin
					state<=17;
					out<=223;
				end
				if(in == 223) begin
					state<=1;
					out<=224;
				end
				if(in == 224) begin
					state<=17;
					out<=225;
				end
				if(in == 225) begin
					state<=1;
					out<=226;
				end
				if(in == 226) begin
					state<=17;
					out<=227;
				end
				if(in == 227) begin
					state<=1;
					out<=228;
				end
				if(in == 228) begin
					state<=17;
					out<=229;
				end
				if(in == 229) begin
					state<=1;
					out<=230;
				end
				if(in == 230) begin
					state<=17;
					out<=231;
				end
				if(in == 231) begin
					state<=1;
					out<=232;
				end
				if(in == 232) begin
					state<=17;
					out<=233;
				end
				if(in == 233) begin
					state<=15;
					out<=234;
				end
				if(in == 234) begin
					state<=17;
					out<=235;
				end
				if(in == 235) begin
					state<=15;
					out<=236;
				end
				if(in == 236) begin
					state<=17;
					out<=237;
				end
				if(in == 237) begin
					state<=15;
					out<=238;
				end
				if(in == 238) begin
					state<=17;
					out<=239;
				end
				if(in == 239) begin
					state<=17;
					out<=240;
				end
				if(in == 240) begin
					state<=17;
					out<=241;
				end
				if(in == 241) begin
					state<=17;
					out<=242;
				end
				if(in == 242) begin
					state<=17;
					out<=243;
				end
				if(in == 243) begin
					state<=17;
					out<=244;
				end
				if(in == 244) begin
					state<=17;
					out<=245;
				end
				if(in == 245) begin
					state<=17;
					out<=246;
				end
				if(in == 246) begin
					state<=17;
					out<=247;
				end
				if(in == 247) begin
					state<=17;
					out<=248;
				end
				if(in == 248) begin
					state<=17;
					out<=249;
				end
				if(in == 249) begin
					state<=17;
					out<=250;
				end
				if(in == 250) begin
					state<=17;
					out<=251;
				end
				if(in == 251) begin
					state<=17;
					out<=252;
				end
				if(in == 252) begin
					state<=17;
					out<=253;
				end
				if(in == 253) begin
					state<=17;
					out<=254;
				end
				if(in == 254) begin
					state<=17;
					out<=255;
				end
				if(in == 255) begin
					state<=17;
					out<=0;
				end
				if(in == 256) begin
					state<=17;
					out<=1;
				end
				if(in == 257) begin
					state<=17;
					out<=2;
				end
				if(in == 258) begin
					state<=17;
					out<=3;
				end
				if(in == 259) begin
					state<=17;
					out<=4;
				end
				if(in == 260) begin
					state<=17;
					out<=5;
				end
				if(in == 261) begin
					state<=17;
					out<=6;
				end
				if(in == 262) begin
					state<=17;
					out<=7;
				end
				if(in == 263) begin
					state<=17;
					out<=8;
				end
				if(in == 264) begin
					state<=17;
					out<=9;
				end
				if(in == 265) begin
					state<=17;
					out<=10;
				end
				if(in == 266) begin
					state<=17;
					out<=11;
				end
				if(in == 267) begin
					state<=17;
					out<=12;
				end
				if(in == 268) begin
					state<=17;
					out<=13;
				end
				if(in == 269) begin
					state<=17;
					out<=14;
				end
				if(in == 270) begin
					state<=17;
					out<=15;
				end
				if(in == 271) begin
					state<=17;
					out<=16;
				end
				if(in == 272) begin
					state<=17;
					out<=17;
				end
				if(in == 273) begin
					state<=17;
					out<=18;
				end
				if(in == 274) begin
					state<=17;
					out<=19;
				end
				if(in == 275) begin
					state<=17;
					out<=20;
				end
				if(in == 276) begin
					state<=17;
					out<=21;
				end
				if(in == 277) begin
					state<=17;
					out<=22;
				end
				if(in == 278) begin
					state<=17;
					out<=23;
				end
				if(in == 279) begin
					state<=17;
					out<=24;
				end
				if(in == 280) begin
					state<=17;
					out<=25;
				end
				if(in == 281) begin
					state<=17;
					out<=26;
				end
				if(in == 282) begin
					state<=17;
					out<=27;
				end
				if(in == 283) begin
					state<=17;
					out<=28;
				end
				if(in == 284) begin
					state<=17;
					out<=29;
				end
				if(in == 285) begin
					state<=15;
					out<=30;
				end
				if(in == 286) begin
					state<=17;
					out<=31;
				end
				if(in == 287) begin
					state<=15;
					out<=32;
				end
				if(in == 288) begin
					state<=17;
					out<=33;
				end
				if(in == 289) begin
					state<=15;
					out<=34;
				end
				if(in == 290) begin
					state<=17;
					out<=35;
				end
				if(in == 291) begin
					state<=17;
					out<=36;
				end
				if(in == 292) begin
					state<=17;
					out<=37;
				end
				if(in == 293) begin
					state<=17;
					out<=38;
				end
				if(in == 294) begin
					state<=17;
					out<=39;
				end
				if(in == 295) begin
					state<=17;
					out<=40;
				end
				if(in == 296) begin
					state<=17;
					out<=41;
				end
				if(in == 297) begin
					state<=17;
					out<=42;
				end
				if(in == 298) begin
					state<=17;
					out<=43;
				end
				if(in == 299) begin
					state<=17;
					out<=44;
				end
				if(in == 300) begin
					state<=17;
					out<=45;
				end
				if(in == 301) begin
					state<=17;
					out<=46;
				end
				if(in == 302) begin
					state<=17;
					out<=47;
				end
				if(in == 303) begin
					state<=17;
					out<=48;
				end
				if(in == 304) begin
					state<=17;
					out<=49;
				end
				if(in == 305) begin
					state<=17;
					out<=50;
				end
				if(in == 306) begin
					state<=17;
					out<=51;
				end
				if(in == 307) begin
					state<=17;
					out<=52;
				end
				if(in == 308) begin
					state<=17;
					out<=53;
				end
				if(in == 309) begin
					state<=17;
					out<=54;
				end
				if(in == 310) begin
					state<=17;
					out<=55;
				end
				if(in == 311) begin
					state<=17;
					out<=56;
				end
				if(in == 312) begin
					state<=17;
					out<=57;
				end
				if(in == 313) begin
					state<=17;
					out<=58;
				end
				if(in == 314) begin
					state<=17;
					out<=59;
				end
				if(in == 315) begin
					state<=17;
					out<=60;
				end
				if(in == 316) begin
					state<=17;
					out<=61;
				end
				if(in == 317) begin
					state<=17;
					out<=62;
				end
				if(in == 318) begin
					state<=17;
					out<=63;
				end
				if(in == 319) begin
					state<=17;
					out<=64;
				end
				if(in == 320) begin
					state<=17;
					out<=65;
				end
				if(in == 321) begin
					state<=17;
					out<=66;
				end
				if(in == 322) begin
					state<=17;
					out<=67;
				end
				if(in == 323) begin
					state<=17;
					out<=68;
				end
				if(in == 324) begin
					state<=17;
					out<=69;
				end
				if(in == 325) begin
					state<=17;
					out<=70;
				end
				if(in == 326) begin
					state<=17;
					out<=71;
				end
				if(in == 327) begin
					state<=17;
					out<=72;
				end
				if(in == 328) begin
					state<=17;
					out<=73;
				end
				if(in == 329) begin
					state<=17;
					out<=74;
				end
				if(in == 330) begin
					state<=17;
					out<=75;
				end
				if(in == 331) begin
					state<=17;
					out<=76;
				end
				if(in == 332) begin
					state<=17;
					out<=77;
				end
				if(in == 333) begin
					state<=17;
					out<=78;
				end
				if(in == 334) begin
					state<=17;
					out<=79;
				end
				if(in == 335) begin
					state<=17;
					out<=80;
				end
				if(in == 336) begin
					state<=17;
					out<=81;
				end
				if(in == 337) begin
					state<=15;
					out<=82;
				end
				if(in == 338) begin
					state<=17;
					out<=83;
				end
				if(in == 339) begin
					state<=15;
					out<=84;
				end
				if(in == 340) begin
					state<=17;
					out<=85;
				end
				if(in == 341) begin
					state<=15;
					out<=86;
				end
				if(in == 342) begin
					state<=17;
					out<=87;
				end
				if(in == 343) begin
					state<=15;
					out<=88;
				end
				if(in == 344) begin
					state<=17;
					out<=89;
				end
				if(in == 345) begin
					state<=15;
					out<=90;
				end
				if(in == 346) begin
					state<=17;
					out<=91;
				end
				if(in == 347) begin
					state<=15;
					out<=92;
				end
				if(in == 348) begin
					state<=17;
					out<=93;
				end
				if(in == 349) begin
					state<=16;
					out<=94;
				end
				if(in == 350) begin
					state<=16;
					out<=95;
				end
				if(in == 351) begin
					state<=16;
					out<=96;
				end
				if(in == 352) begin
					state<=16;
					out<=97;
				end
				if(in == 353) begin
					state<=16;
					out<=98;
				end
				if(in == 354) begin
					state<=16;
					out<=99;
				end
				if(in == 355) begin
					state<=16;
					out<=100;
				end
				if(in == 356) begin
					state<=16;
					out<=101;
				end
				if(in == 357) begin
					state<=16;
					out<=102;
				end
				if(in == 358) begin
					state<=16;
					out<=103;
				end
				if(in == 359) begin
					state<=16;
					out<=104;
				end
				if(in == 360) begin
					state<=16;
					out<=105;
				end
				if(in == 361) begin
					state<=16;
					out<=106;
				end
				if(in == 362) begin
					state<=16;
					out<=107;
				end
				if(in == 363) begin
					state<=16;
					out<=108;
				end
				if(in == 364) begin
					state<=16;
					out<=109;
				end
				if(in == 365) begin
					state<=16;
					out<=110;
				end
				if(in == 366) begin
					state<=16;
					out<=111;
				end
				if(in == 367) begin
					state<=16;
					out<=112;
				end
				if(in == 368) begin
					state<=16;
					out<=113;
				end
				if(in == 369) begin
					state<=16;
					out<=114;
				end
				if(in == 370) begin
					state<=16;
					out<=115;
				end
				if(in == 371) begin
					state<=16;
					out<=116;
				end
				if(in == 372) begin
					state<=16;
					out<=117;
				end
				if(in == 373) begin
					state<=16;
					out<=118;
				end
				if(in == 374) begin
					state<=16;
					out<=119;
				end
				if(in == 375) begin
					state<=16;
					out<=120;
				end
				if(in == 376) begin
					state<=16;
					out<=121;
				end
				if(in == 377) begin
					state<=16;
					out<=122;
				end
				if(in == 378) begin
					state<=16;
					out<=123;
				end
				if(in == 379) begin
					state<=16;
					out<=124;
				end
				if(in == 380) begin
					state<=16;
					out<=125;
				end
				if(in == 381) begin
					state<=16;
					out<=126;
				end
				if(in == 382) begin
					state<=16;
					out<=127;
				end
				if(in == 383) begin
					state<=16;
					out<=128;
				end
				if(in == 384) begin
					state<=16;
					out<=129;
				end
				if(in == 385) begin
					state<=16;
					out<=130;
				end
				if(in == 386) begin
					state<=16;
					out<=131;
				end
				if(in == 387) begin
					state<=16;
					out<=132;
				end
				if(in == 388) begin
					state<=16;
					out<=133;
				end
				if(in == 389) begin
					state<=16;
					out<=134;
				end
				if(in == 390) begin
					state<=16;
					out<=135;
				end
				if(in == 391) begin
					state<=16;
					out<=136;
				end
				if(in == 392) begin
					state<=16;
					out<=137;
				end
				if(in == 393) begin
					state<=16;
					out<=138;
				end
				if(in == 394) begin
					state<=16;
					out<=139;
				end
				if(in == 395) begin
					state<=16;
					out<=140;
				end
				if(in == 396) begin
					state<=16;
					out<=141;
				end
				if(in == 397) begin
					state<=16;
					out<=142;
				end
				if(in == 398) begin
					state<=16;
					out<=143;
				end
				if(in == 399) begin
					state<=16;
					out<=144;
				end
				if(in == 400) begin
					state<=16;
					out<=145;
				end
				if(in == 401) begin
					state<=16;
					out<=146;
				end
				if(in == 402) begin
					state<=16;
					out<=147;
				end
				if(in == 403) begin
					state<=16;
					out<=148;
				end
				if(in == 404) begin
					state<=16;
					out<=149;
				end
				if(in == 405) begin
					state<=16;
					out<=150;
				end
				if(in == 406) begin
					state<=16;
					out<=151;
				end
				if(in == 407) begin
					state<=16;
					out<=152;
				end
				if(in == 408) begin
					state<=16;
					out<=153;
				end
				if(in == 409) begin
					state<=16;
					out<=154;
				end
				if(in == 410) begin
					state<=16;
					out<=155;
				end
				if(in == 411) begin
					state<=16;
					out<=156;
				end
				if(in == 412) begin
					state<=16;
					out<=157;
				end
				if(in == 413) begin
					state<=16;
					out<=158;
				end
				if(in == 414) begin
					state<=16;
					out<=159;
				end
				if(in == 415) begin
					state<=16;
					out<=160;
				end
				if(in == 416) begin
					state<=16;
					out<=161;
				end
				if(in == 417) begin
					state<=16;
					out<=162;
				end
				if(in == 418) begin
					state<=16;
					out<=163;
				end
				if(in == 419) begin
					state<=16;
					out<=164;
				end
				if(in == 420) begin
					state<=16;
					out<=165;
				end
				if(in == 421) begin
					state<=16;
					out<=166;
				end
				if(in == 422) begin
					state<=16;
					out<=167;
				end
				if(in == 423) begin
					state<=16;
					out<=168;
				end
				if(in == 424) begin
					state<=16;
					out<=169;
				end
				if(in == 425) begin
					state<=16;
					out<=170;
				end
				if(in == 426) begin
					state<=16;
					out<=171;
				end
				if(in == 427) begin
					state<=16;
					out<=172;
				end
				if(in == 428) begin
					state<=16;
					out<=173;
				end
				if(in == 429) begin
					state<=16;
					out<=174;
				end
				if(in == 430) begin
					state<=16;
					out<=175;
				end
				if(in == 431) begin
					state<=16;
					out<=176;
				end
				if(in == 432) begin
					state<=16;
					out<=177;
				end
				if(in == 433) begin
					state<=16;
					out<=178;
				end
				if(in == 434) begin
					state<=16;
					out<=179;
				end
				if(in == 435) begin
					state<=16;
					out<=180;
				end
				if(in == 436) begin
					state<=16;
					out<=181;
				end
				if(in == 437) begin
					state<=16;
					out<=182;
				end
				if(in == 438) begin
					state<=16;
					out<=183;
				end
				if(in == 439) begin
					state<=16;
					out<=184;
				end
				if(in == 440) begin
					state<=16;
					out<=185;
				end
				if(in == 441) begin
					state<=16;
					out<=186;
				end
				if(in == 442) begin
					state<=16;
					out<=187;
				end
				if(in == 443) begin
					state<=16;
					out<=188;
				end
				if(in == 444) begin
					state<=16;
					out<=189;
				end
				if(in == 445) begin
					state<=16;
					out<=190;
				end
				if(in == 446) begin
					state<=16;
					out<=191;
				end
				if(in == 447) begin
					state<=16;
					out<=192;
				end
				if(in == 448) begin
					state<=16;
					out<=193;
				end
				if(in == 449) begin
					state<=16;
					out<=194;
				end
				if(in == 450) begin
					state<=16;
					out<=195;
				end
				if(in == 451) begin
					state<=16;
					out<=196;
				end
				if(in == 452) begin
					state<=16;
					out<=197;
				end
				if(in == 453) begin
					state<=16;
					out<=198;
				end
				if(in == 454) begin
					state<=16;
					out<=199;
				end
				if(in == 455) begin
					state<=16;
					out<=200;
				end
				if(in == 456) begin
					state<=16;
					out<=201;
				end
				if(in == 457) begin
					state<=16;
					out<=202;
				end
				if(in == 458) begin
					state<=16;
					out<=203;
				end
				if(in == 459) begin
					state<=16;
					out<=204;
				end
				if(in == 460) begin
					state<=16;
					out<=205;
				end
				if(in == 461) begin
					state<=16;
					out<=206;
				end
				if(in == 462) begin
					state<=16;
					out<=207;
				end
				if(in == 463) begin
					state<=16;
					out<=208;
				end
				if(in == 464) begin
					state<=16;
					out<=209;
				end
				if(in == 465) begin
					state<=1;
					out<=210;
				end
				if(in == 466) begin
					state<=17;
					out<=211;
				end
				if(in == 467) begin
					state<=1;
					out<=212;
				end
				if(in == 468) begin
					state<=17;
					out<=213;
				end
				if(in == 469) begin
					state<=1;
					out<=214;
				end
				if(in == 470) begin
					state<=17;
					out<=215;
				end
				if(in == 471) begin
					state<=17;
					out<=216;
				end
				if(in == 472) begin
					state<=17;
					out<=217;
				end
				if(in == 473) begin
					state<=17;
					out<=218;
				end
				if(in == 474) begin
					state<=17;
					out<=219;
				end
				if(in == 475) begin
					state<=17;
					out<=220;
				end
				if(in == 476) begin
					state<=17;
					out<=221;
				end
				if(in == 477) begin
					state<=17;
					out<=222;
				end
				if(in == 478) begin
					state<=17;
					out<=223;
				end
				if(in == 479) begin
					state<=17;
					out<=224;
				end
				if(in == 480) begin
					state<=17;
					out<=225;
				end
				if(in == 481) begin
					state<=17;
					out<=226;
				end
				if(in == 482) begin
					state<=17;
					out<=227;
				end
				if(in == 483) begin
					state<=17;
					out<=228;
				end
				if(in == 484) begin
					state<=17;
					out<=229;
				end
				if(in == 485) begin
					state<=17;
					out<=230;
				end
				if(in == 486) begin
					state<=17;
					out<=231;
				end
				if(in == 487) begin
					state<=17;
					out<=232;
				end
				if(in == 488) begin
					state<=17;
					out<=233;
				end
				if(in == 489) begin
					state<=17;
					out<=234;
				end
				if(in == 490) begin
					state<=17;
					out<=235;
				end
				if(in == 491) begin
					state<=17;
					out<=236;
				end
				if(in == 492) begin
					state<=17;
					out<=237;
				end
				if(in == 493) begin
					state<=17;
					out<=238;
				end
				if(in == 494) begin
					state<=17;
					out<=239;
				end
				if(in == 495) begin
					state<=17;
					out<=240;
				end
				if(in == 496) begin
					state<=17;
					out<=241;
				end
				if(in == 497) begin
					state<=17;
					out<=242;
				end
				if(in == 498) begin
					state<=17;
					out<=243;
				end
				if(in == 499) begin
					state<=17;
					out<=244;
				end
				if(in == 500) begin
					state<=17;
					out<=245;
				end
				if(in == 501) begin
					state<=17;
					out<=246;
				end
				if(in == 502) begin
					state<=17;
					out<=247;
				end
				if(in == 503) begin
					state<=17;
					out<=248;
				end
				if(in == 504) begin
					state<=17;
					out<=249;
				end
				if(in == 505) begin
					state<=17;
					out<=250;
				end
				if(in == 506) begin
					state<=17;
					out<=251;
				end
				if(in == 507) begin
					state<=17;
					out<=252;
				end
				if(in == 508) begin
					state<=17;
					out<=253;
				end
				if(in == 509) begin
					state<=17;
					out<=254;
				end
				if(in == 510) begin
					state<=17;
					out<=255;
				end
				if(in == 511) begin
					state<=17;
					out<=0;
				end
				if(in == 512) begin
					state<=17;
					out<=1;
				end
				if(in == 513) begin
					state<=17;
					out<=2;
				end
				if(in == 514) begin
					state<=17;
					out<=3;
				end
				if(in == 515) begin
					state<=17;
					out<=4;
				end
				if(in == 516) begin
					state<=17;
					out<=5;
				end
				if(in == 517) begin
					state<=1;
					out<=6;
				end
				if(in == 518) begin
					state<=17;
					out<=7;
				end
				if(in == 519) begin
					state<=1;
					out<=8;
				end
				if(in == 520) begin
					state<=17;
					out<=9;
				end
				if(in == 521) begin
					state<=1;
					out<=10;
				end
				if(in == 522) begin
					state<=17;
					out<=11;
				end
				if(in == 523) begin
					state<=17;
					out<=12;
				end
				if(in == 524) begin
					state<=17;
					out<=13;
				end
				if(in == 525) begin
					state<=17;
					out<=14;
				end
				if(in == 526) begin
					state<=17;
					out<=15;
				end
				if(in == 527) begin
					state<=17;
					out<=16;
				end
				if(in == 528) begin
					state<=17;
					out<=17;
				end
				if(in == 529) begin
					state<=17;
					out<=18;
				end
				if(in == 530) begin
					state<=17;
					out<=19;
				end
				if(in == 531) begin
					state<=17;
					out<=20;
				end
				if(in == 532) begin
					state<=17;
					out<=21;
				end
				if(in == 533) begin
					state<=17;
					out<=22;
				end
				if(in == 534) begin
					state<=17;
					out<=23;
				end
				if(in == 535) begin
					state<=17;
					out<=24;
				end
				if(in == 536) begin
					state<=17;
					out<=25;
				end
				if(in == 537) begin
					state<=17;
					out<=26;
				end
				if(in == 538) begin
					state<=17;
					out<=27;
				end
				if(in == 539) begin
					state<=17;
					out<=28;
				end
				if(in == 540) begin
					state<=17;
					out<=29;
				end
				if(in == 541) begin
					state<=17;
					out<=30;
				end
				if(in == 542) begin
					state<=17;
					out<=31;
				end
				if(in == 543) begin
					state<=17;
					out<=32;
				end
				if(in == 544) begin
					state<=17;
					out<=33;
				end
				if(in == 545) begin
					state<=17;
					out<=34;
				end
				if(in == 546) begin
					state<=17;
					out<=35;
				end
				if(in == 547) begin
					state<=17;
					out<=36;
				end
				if(in == 548) begin
					state<=17;
					out<=37;
				end
				if(in == 549) begin
					state<=17;
					out<=38;
				end
				if(in == 550) begin
					state<=17;
					out<=39;
				end
				if(in == 551) begin
					state<=17;
					out<=40;
				end
				if(in == 552) begin
					state<=17;
					out<=41;
				end
				if(in == 553) begin
					state<=17;
					out<=42;
				end
				if(in == 554) begin
					state<=17;
					out<=43;
				end
				if(in == 555) begin
					state<=17;
					out<=44;
				end
				if(in == 556) begin
					state<=17;
					out<=45;
				end
				if(in == 557) begin
					state<=17;
					out<=46;
				end
				if(in == 558) begin
					state<=17;
					out<=47;
				end
				if(in == 559) begin
					state<=17;
					out<=48;
				end
				if(in == 560) begin
					state<=17;
					out<=49;
				end
				if(in == 561) begin
					state<=17;
					out<=50;
				end
				if(in == 562) begin
					state<=17;
					out<=51;
				end
				if(in == 563) begin
					state<=17;
					out<=52;
				end
				if(in == 564) begin
					state<=17;
					out<=53;
				end
				if(in == 565) begin
					state<=17;
					out<=54;
				end
				if(in == 566) begin
					state<=17;
					out<=55;
				end
				if(in == 567) begin
					state<=17;
					out<=56;
				end
				if(in == 568) begin
					state<=17;
					out<=57;
				end
				if(in == 569) begin
					state<=1;
					out<=58;
				end
				if(in == 570) begin
					state<=17;
					out<=59;
				end
				if(in == 571) begin
					state<=1;
					out<=60;
				end
				if(in == 572) begin
					state<=17;
					out<=61;
				end
				if(in == 573) begin
					state<=1;
					out<=62;
				end
				if(in == 574) begin
					state<=17;
					out<=63;
				end
				if(in == 575) begin
					state<=1;
					out<=64;
				end
				if(in == 576) begin
					state<=17;
					out<=65;
				end
				if(in == 577) begin
					state<=1;
					out<=66;
				end
				if(in == 578) begin
					state<=17;
					out<=67;
				end
				if(in == 579) begin
					state<=1;
					out<=68;
				end
				if(in == 580) begin
					state<=17;
					out<=69;
				end
				if(in == 581) begin
					state<=1;
					out<=70;
				end
				if(in == 582) begin
					state<=17;
					out<=71;
				end
				if(in == 583) begin
					state<=1;
					out<=72;
				end
				if(in == 584) begin
					state<=17;
					out<=73;
				end
				if(in == 585) begin
					state<=1;
					out<=74;
				end
				if(in == 586) begin
					state<=17;
					out<=75;
				end
				if(in == 587) begin
					state<=17;
					out<=76;
				end
				if(in == 588) begin
					state<=17;
					out<=77;
				end
				if(in == 589) begin
					state<=17;
					out<=78;
				end
				if(in == 590) begin
					state<=17;
					out<=79;
				end
				if(in == 591) begin
					state<=17;
					out<=80;
				end
				if(in == 592) begin
					state<=17;
					out<=81;
				end
				if(in == 593) begin
					state<=17;
					out<=82;
				end
				if(in == 594) begin
					state<=17;
					out<=83;
				end
				if(in == 595) begin
					state<=17;
					out<=84;
				end
				if(in == 596) begin
					state<=17;
					out<=85;
				end
				if(in == 597) begin
					state<=17;
					out<=86;
				end
				if(in == 598) begin
					state<=17;
					out<=87;
				end
				if(in == 599) begin
					state<=17;
					out<=88;
				end
				if(in == 600) begin
					state<=17;
					out<=89;
				end
				if(in == 601) begin
					state<=17;
					out<=90;
				end
				if(in == 602) begin
					state<=17;
					out<=91;
				end
				if(in == 603) begin
					state<=17;
					out<=92;
				end
				if(in == 604) begin
					state<=17;
					out<=93;
				end
				if(in == 605) begin
					state<=17;
					out<=94;
				end
				if(in == 606) begin
					state<=17;
					out<=95;
				end
				if(in == 607) begin
					state<=17;
					out<=96;
				end
				if(in == 608) begin
					state<=17;
					out<=97;
				end
				if(in == 609) begin
					state<=17;
					out<=98;
				end
				if(in == 610) begin
					state<=17;
					out<=99;
				end
				if(in == 611) begin
					state<=17;
					out<=100;
				end
				if(in == 612) begin
					state<=17;
					out<=101;
				end
				if(in == 613) begin
					state<=17;
					out<=102;
				end
				if(in == 614) begin
					state<=17;
					out<=103;
				end
				if(in == 615) begin
					state<=17;
					out<=104;
				end
				if(in == 616) begin
					state<=17;
					out<=105;
				end
				if(in == 617) begin
					state<=17;
					out<=106;
				end
				if(in == 618) begin
					state<=17;
					out<=107;
				end
				if(in == 619) begin
					state<=17;
					out<=108;
				end
				if(in == 620) begin
					state<=17;
					out<=109;
				end
				if(in == 621) begin
					state<=17;
					out<=110;
				end
				if(in == 622) begin
					state<=17;
					out<=111;
				end
				if(in == 623) begin
					state<=17;
					out<=112;
				end
				if(in == 624) begin
					state<=17;
					out<=113;
				end
				if(in == 625) begin
					state<=17;
					out<=114;
				end
				if(in == 626) begin
					state<=17;
					out<=115;
				end
				if(in == 627) begin
					state<=17;
					out<=116;
				end
				if(in == 628) begin
					state<=17;
					out<=117;
				end
				if(in == 629) begin
					state<=17;
					out<=118;
				end
				if(in == 630) begin
					state<=17;
					out<=119;
				end
				if(in == 631) begin
					state<=17;
					out<=120;
				end
				if(in == 632) begin
					state<=17;
					out<=121;
				end
				if(in == 633) begin
					state<=1;
					out<=122;
				end
				if(in == 634) begin
					state<=17;
					out<=123;
				end
				if(in == 635) begin
					state<=1;
					out<=124;
				end
				if(in == 636) begin
					state<=17;
					out<=125;
				end
				if(in == 637) begin
					state<=1;
					out<=126;
				end
				if(in == 638) begin
					state<=17;
					out<=127;
				end
				if(in == 639) begin
					state<=17;
					out<=128;
				end
				if(in == 640) begin
					state<=17;
					out<=129;
				end
				if(in == 641) begin
					state<=17;
					out<=130;
				end
				if(in == 642) begin
					state<=17;
					out<=131;
				end
				if(in == 643) begin
					state<=17;
					out<=132;
				end
				if(in == 644) begin
					state<=17;
					out<=133;
				end
				if(in == 645) begin
					state<=17;
					out<=134;
				end
				if(in == 646) begin
					state<=17;
					out<=135;
				end
				if(in == 647) begin
					state<=17;
					out<=136;
				end
				if(in == 648) begin
					state<=17;
					out<=137;
				end
				if(in == 649) begin
					state<=17;
					out<=138;
				end
				if(in == 650) begin
					state<=17;
					out<=139;
				end
				if(in == 651) begin
					state<=17;
					out<=140;
				end
				if(in == 652) begin
					state<=17;
					out<=141;
				end
				if(in == 653) begin
					state<=17;
					out<=142;
				end
				if(in == 654) begin
					state<=17;
					out<=143;
				end
				if(in == 655) begin
					state<=17;
					out<=144;
				end
				if(in == 656) begin
					state<=17;
					out<=145;
				end
				if(in == 657) begin
					state<=17;
					out<=146;
				end
				if(in == 658) begin
					state<=17;
					out<=147;
				end
				if(in == 659) begin
					state<=17;
					out<=148;
				end
				if(in == 660) begin
					state<=17;
					out<=149;
				end
				if(in == 661) begin
					state<=17;
					out<=150;
				end
				if(in == 662) begin
					state<=17;
					out<=151;
				end
				if(in == 663) begin
					state<=17;
					out<=152;
				end
				if(in == 664) begin
					state<=17;
					out<=153;
				end
				if(in == 665) begin
					state<=17;
					out<=154;
				end
				if(in == 666) begin
					state<=17;
					out<=155;
				end
				if(in == 667) begin
					state<=17;
					out<=156;
				end
				if(in == 668) begin
					state<=17;
					out<=157;
				end
				if(in == 669) begin
					state<=17;
					out<=158;
				end
				if(in == 670) begin
					state<=17;
					out<=159;
				end
				if(in == 671) begin
					state<=17;
					out<=160;
				end
				if(in == 672) begin
					state<=17;
					out<=161;
				end
				if(in == 673) begin
					state<=17;
					out<=162;
				end
				if(in == 674) begin
					state<=17;
					out<=163;
				end
				if(in == 675) begin
					state<=17;
					out<=164;
				end
				if(in == 676) begin
					state<=17;
					out<=165;
				end
				if(in == 677) begin
					state<=17;
					out<=166;
				end
				if(in == 678) begin
					state<=17;
					out<=167;
				end
				if(in == 679) begin
					state<=17;
					out<=168;
				end
				if(in == 680) begin
					state<=17;
					out<=169;
				end
				if(in == 681) begin
					state<=17;
					out<=170;
				end
				if(in == 682) begin
					state<=17;
					out<=171;
				end
				if(in == 683) begin
					state<=17;
					out<=172;
				end
				if(in == 684) begin
					state<=17;
					out<=173;
				end
				if(in == 685) begin
					state<=1;
					out<=174;
				end
				if(in == 686) begin
					state<=17;
					out<=175;
				end
				if(in == 687) begin
					state<=1;
					out<=176;
				end
				if(in == 688) begin
					state<=17;
					out<=177;
				end
				if(in == 689) begin
					state<=1;
					out<=178;
				end
				if(in == 690) begin
					state<=17;
					out<=179;
				end
				if(in == 691) begin
					state<=1;
					out<=180;
				end
				if(in == 692) begin
					state<=17;
					out<=181;
				end
				if(in == 693) begin
					state<=1;
					out<=182;
				end
				if(in == 694) begin
					state<=17;
					out<=183;
				end
				if(in == 695) begin
					state<=1;
					out<=184;
				end
				if(in == 696) begin
					state<=17;
					out<=185;
				end
				if(in == 697) begin
					state<=15;
					out<=186;
				end
				if(in == 698) begin
					state<=17;
					out<=187;
				end
				if(in == 699) begin
					state<=15;
					out<=188;
				end
				if(in == 700) begin
					state<=17;
					out<=189;
				end
				if(in == 701) begin
					state<=15;
					out<=190;
				end
				if(in == 702) begin
					state<=17;
					out<=191;
				end
				if(in == 703) begin
					state<=17;
					out<=192;
				end
				if(in == 704) begin
					state<=17;
					out<=193;
				end
				if(in == 705) begin
					state<=17;
					out<=194;
				end
				if(in == 706) begin
					state<=17;
					out<=195;
				end
				if(in == 707) begin
					state<=17;
					out<=196;
				end
				if(in == 708) begin
					state<=17;
					out<=197;
				end
				if(in == 709) begin
					state<=17;
					out<=198;
				end
				if(in == 710) begin
					state<=17;
					out<=199;
				end
				if(in == 711) begin
					state<=17;
					out<=200;
				end
				if(in == 712) begin
					state<=17;
					out<=201;
				end
				if(in == 713) begin
					state<=17;
					out<=202;
				end
				if(in == 714) begin
					state<=17;
					out<=203;
				end
				if(in == 715) begin
					state<=17;
					out<=204;
				end
				if(in == 716) begin
					state<=17;
					out<=205;
				end
				if(in == 717) begin
					state<=17;
					out<=206;
				end
				if(in == 718) begin
					state<=17;
					out<=207;
				end
				if(in == 719) begin
					state<=17;
					out<=208;
				end
				if(in == 720) begin
					state<=17;
					out<=209;
				end
				if(in == 721) begin
					state<=17;
					out<=210;
				end
				if(in == 722) begin
					state<=17;
					out<=211;
				end
				if(in == 723) begin
					state<=17;
					out<=212;
				end
				if(in == 724) begin
					state<=17;
					out<=213;
				end
				if(in == 725) begin
					state<=17;
					out<=214;
				end
				if(in == 726) begin
					state<=17;
					out<=215;
				end
				if(in == 727) begin
					state<=17;
					out<=216;
				end
				if(in == 728) begin
					state<=17;
					out<=217;
				end
				if(in == 729) begin
					state<=17;
					out<=218;
				end
				if(in == 730) begin
					state<=17;
					out<=219;
				end
				if(in == 731) begin
					state<=17;
					out<=220;
				end
				if(in == 732) begin
					state<=17;
					out<=221;
				end
				if(in == 733) begin
					state<=17;
					out<=222;
				end
				if(in == 734) begin
					state<=17;
					out<=223;
				end
				if(in == 735) begin
					state<=17;
					out<=224;
				end
				if(in == 736) begin
					state<=17;
					out<=225;
				end
				if(in == 737) begin
					state<=17;
					out<=226;
				end
				if(in == 738) begin
					state<=17;
					out<=227;
				end
				if(in == 739) begin
					state<=17;
					out<=228;
				end
				if(in == 740) begin
					state<=17;
					out<=229;
				end
				if(in == 741) begin
					state<=17;
					out<=230;
				end
				if(in == 742) begin
					state<=17;
					out<=231;
				end
				if(in == 743) begin
					state<=17;
					out<=232;
				end
				if(in == 744) begin
					state<=17;
					out<=233;
				end
				if(in == 745) begin
					state<=17;
					out<=234;
				end
				if(in == 746) begin
					state<=17;
					out<=235;
				end
				if(in == 747) begin
					state<=17;
					out<=236;
				end
				if(in == 748) begin
					state<=17;
					out<=237;
				end
				if(in == 749) begin
					state<=15;
					out<=238;
				end
				if(in == 750) begin
					state<=17;
					out<=239;
				end
				if(in == 751) begin
					state<=15;
					out<=240;
				end
				if(in == 752) begin
					state<=17;
					out<=241;
				end
				if(in == 753) begin
					state<=15;
					out<=242;
				end
				if(in == 754) begin
					state<=17;
					out<=243;
				end
				if(in == 755) begin
					state<=17;
					out<=244;
				end
				if(in == 756) begin
					state<=17;
					out<=245;
				end
				if(in == 757) begin
					state<=17;
					out<=246;
				end
				if(in == 758) begin
					state<=17;
					out<=247;
				end
				if(in == 759) begin
					state<=17;
					out<=248;
				end
				if(in == 760) begin
					state<=17;
					out<=249;
				end
				if(in == 761) begin
					state<=17;
					out<=250;
				end
				if(in == 762) begin
					state<=17;
					out<=251;
				end
				if(in == 763) begin
					state<=17;
					out<=252;
				end
				if(in == 764) begin
					state<=17;
					out<=253;
				end
				if(in == 765) begin
					state<=17;
					out<=254;
				end
				if(in == 766) begin
					state<=17;
					out<=255;
				end
				if(in == 767) begin
					state<=17;
					out<=0;
				end
				if(in == 768) begin
					state<=17;
					out<=1;
				end
				if(in == 769) begin
					state<=17;
					out<=2;
				end
				if(in == 770) begin
					state<=17;
					out<=3;
				end
				if(in == 771) begin
					state<=17;
					out<=4;
				end
				if(in == 772) begin
					state<=17;
					out<=5;
				end
				if(in == 773) begin
					state<=17;
					out<=6;
				end
				if(in == 774) begin
					state<=17;
					out<=7;
				end
				if(in == 775) begin
					state<=17;
					out<=8;
				end
				if(in == 776) begin
					state<=17;
					out<=9;
				end
				if(in == 777) begin
					state<=17;
					out<=10;
				end
				if(in == 778) begin
					state<=17;
					out<=11;
				end
				if(in == 779) begin
					state<=17;
					out<=12;
				end
				if(in == 780) begin
					state<=17;
					out<=13;
				end
				if(in == 781) begin
					state<=17;
					out<=14;
				end
				if(in == 782) begin
					state<=17;
					out<=15;
				end
				if(in == 783) begin
					state<=17;
					out<=16;
				end
				if(in == 784) begin
					state<=17;
					out<=17;
				end
				if(in == 785) begin
					state<=17;
					out<=18;
				end
				if(in == 786) begin
					state<=17;
					out<=19;
				end
				if(in == 787) begin
					state<=17;
					out<=20;
				end
				if(in == 788) begin
					state<=17;
					out<=21;
				end
				if(in == 789) begin
					state<=17;
					out<=22;
				end
				if(in == 790) begin
					state<=17;
					out<=23;
				end
				if(in == 791) begin
					state<=17;
					out<=24;
				end
				if(in == 792) begin
					state<=17;
					out<=25;
				end
				if(in == 793) begin
					state<=17;
					out<=26;
				end
				if(in == 794) begin
					state<=17;
					out<=27;
				end
				if(in == 795) begin
					state<=17;
					out<=28;
				end
				if(in == 796) begin
					state<=17;
					out<=29;
				end
				if(in == 797) begin
					state<=17;
					out<=30;
				end
				if(in == 798) begin
					state<=17;
					out<=31;
				end
				if(in == 799) begin
					state<=17;
					out<=32;
				end
				if(in == 800) begin
					state<=17;
					out<=33;
				end
				if(in == 801) begin
					state<=15;
					out<=34;
				end
				if(in == 802) begin
					state<=17;
					out<=35;
				end
				if(in == 803) begin
					state<=15;
					out<=36;
				end
				if(in == 804) begin
					state<=17;
					out<=37;
				end
				if(in == 805) begin
					state<=15;
					out<=38;
				end
				if(in == 806) begin
					state<=17;
					out<=39;
				end
				if(in == 807) begin
					state<=15;
					out<=40;
				end
				if(in == 808) begin
					state<=17;
					out<=41;
				end
				if(in == 809) begin
					state<=15;
					out<=42;
				end
				if(in == 810) begin
					state<=17;
					out<=43;
				end
				if(in == 811) begin
					state<=15;
					out<=44;
				end
				if(in == 812) begin
					state<=17;
					out<=45;
				end
				if(in == 813) begin
					state<=16;
					out<=46;
				end
				if(in == 814) begin
					state<=16;
					out<=47;
				end
				if(in == 815) begin
					state<=16;
					out<=48;
				end
				if(in == 816) begin
					state<=16;
					out<=49;
				end
				if(in == 817) begin
					state<=16;
					out<=50;
				end
				if(in == 818) begin
					state<=16;
					out<=51;
				end
				if(in == 819) begin
					state<=16;
					out<=52;
				end
				if(in == 820) begin
					state<=16;
					out<=53;
				end
				if(in == 821) begin
					state<=16;
					out<=54;
				end
				if(in == 822) begin
					state<=16;
					out<=55;
				end
				if(in == 823) begin
					state<=16;
					out<=56;
				end
				if(in == 824) begin
					state<=16;
					out<=57;
				end
				if(in == 825) begin
					state<=16;
					out<=58;
				end
				if(in == 826) begin
					state<=16;
					out<=59;
				end
				if(in == 827) begin
					state<=16;
					out<=60;
				end
				if(in == 828) begin
					state<=16;
					out<=61;
				end
				if(in == 829) begin
					state<=16;
					out<=62;
				end
				if(in == 830) begin
					state<=16;
					out<=63;
				end
				if(in == 831) begin
					state<=16;
					out<=64;
				end
				if(in == 832) begin
					state<=16;
					out<=65;
				end
				if(in == 833) begin
					state<=16;
					out<=66;
				end
				if(in == 834) begin
					state<=16;
					out<=67;
				end
				if(in == 835) begin
					state<=16;
					out<=68;
				end
				if(in == 836) begin
					state<=16;
					out<=69;
				end
				if(in == 837) begin
					state<=16;
					out<=70;
				end
				if(in == 838) begin
					state<=16;
					out<=71;
				end
				if(in == 839) begin
					state<=16;
					out<=72;
				end
				if(in == 840) begin
					state<=16;
					out<=73;
				end
				if(in == 841) begin
					state<=16;
					out<=74;
				end
				if(in == 842) begin
					state<=16;
					out<=75;
				end
				if(in == 843) begin
					state<=16;
					out<=76;
				end
				if(in == 844) begin
					state<=16;
					out<=77;
				end
				if(in == 845) begin
					state<=16;
					out<=78;
				end
				if(in == 846) begin
					state<=16;
					out<=79;
				end
				if(in == 847) begin
					state<=16;
					out<=80;
				end
				if(in == 848) begin
					state<=16;
					out<=81;
				end
				if(in == 849) begin
					state<=16;
					out<=82;
				end
				if(in == 850) begin
					state<=16;
					out<=83;
				end
				if(in == 851) begin
					state<=16;
					out<=84;
				end
				if(in == 852) begin
					state<=16;
					out<=85;
				end
				if(in == 853) begin
					state<=16;
					out<=86;
				end
				if(in == 854) begin
					state<=16;
					out<=87;
				end
				if(in == 855) begin
					state<=16;
					out<=88;
				end
				if(in == 856) begin
					state<=16;
					out<=89;
				end
				if(in == 857) begin
					state<=16;
					out<=90;
				end
				if(in == 858) begin
					state<=16;
					out<=91;
				end
				if(in == 859) begin
					state<=16;
					out<=92;
				end
				if(in == 860) begin
					state<=16;
					out<=93;
				end
				if(in == 861) begin
					state<=16;
					out<=94;
				end
				if(in == 862) begin
					state<=16;
					out<=95;
				end
				if(in == 863) begin
					state<=16;
					out<=96;
				end
				if(in == 864) begin
					state<=16;
					out<=97;
				end
				if(in == 865) begin
					state<=16;
					out<=98;
				end
				if(in == 866) begin
					state<=16;
					out<=99;
				end
				if(in == 867) begin
					state<=16;
					out<=100;
				end
				if(in == 868) begin
					state<=16;
					out<=101;
				end
				if(in == 869) begin
					state<=16;
					out<=102;
				end
				if(in == 870) begin
					state<=16;
					out<=103;
				end
				if(in == 871) begin
					state<=16;
					out<=104;
				end
				if(in == 872) begin
					state<=16;
					out<=105;
				end
				if(in == 873) begin
					state<=16;
					out<=106;
				end
				if(in == 874) begin
					state<=16;
					out<=107;
				end
				if(in == 875) begin
					state<=16;
					out<=108;
				end
				if(in == 876) begin
					state<=16;
					out<=109;
				end
				if(in == 877) begin
					state<=16;
					out<=110;
				end
				if(in == 878) begin
					state<=16;
					out<=111;
				end
				if(in == 879) begin
					state<=16;
					out<=112;
				end
				if(in == 880) begin
					state<=16;
					out<=113;
				end
				if(in == 881) begin
					state<=16;
					out<=114;
				end
				if(in == 882) begin
					state<=16;
					out<=115;
				end
				if(in == 883) begin
					state<=16;
					out<=116;
				end
				if(in == 884) begin
					state<=16;
					out<=117;
				end
				if(in == 885) begin
					state<=16;
					out<=118;
				end
				if(in == 886) begin
					state<=16;
					out<=119;
				end
				if(in == 887) begin
					state<=16;
					out<=120;
				end
				if(in == 888) begin
					state<=16;
					out<=121;
				end
				if(in == 889) begin
					state<=16;
					out<=122;
				end
				if(in == 890) begin
					state<=16;
					out<=123;
				end
				if(in == 891) begin
					state<=16;
					out<=124;
				end
				if(in == 892) begin
					state<=16;
					out<=125;
				end
				if(in == 893) begin
					state<=16;
					out<=126;
				end
				if(in == 894) begin
					state<=16;
					out<=127;
				end
				if(in == 895) begin
					state<=16;
					out<=128;
				end
				if(in == 896) begin
					state<=16;
					out<=129;
				end
				if(in == 897) begin
					state<=16;
					out<=130;
				end
				if(in == 898) begin
					state<=16;
					out<=131;
				end
				if(in == 899) begin
					state<=16;
					out<=132;
				end
				if(in == 900) begin
					state<=16;
					out<=133;
				end
				if(in == 901) begin
					state<=16;
					out<=134;
				end
				if(in == 902) begin
					state<=16;
					out<=135;
				end
				if(in == 903) begin
					state<=16;
					out<=136;
				end
				if(in == 904) begin
					state<=16;
					out<=137;
				end
				if(in == 905) begin
					state<=16;
					out<=138;
				end
				if(in == 906) begin
					state<=16;
					out<=139;
				end
				if(in == 907) begin
					state<=16;
					out<=140;
				end
				if(in == 908) begin
					state<=16;
					out<=141;
				end
				if(in == 909) begin
					state<=16;
					out<=142;
				end
				if(in == 910) begin
					state<=16;
					out<=143;
				end
				if(in == 911) begin
					state<=16;
					out<=144;
				end
				if(in == 912) begin
					state<=16;
					out<=145;
				end
				if(in == 913) begin
					state<=16;
					out<=146;
				end
				if(in == 914) begin
					state<=16;
					out<=147;
				end
				if(in == 915) begin
					state<=16;
					out<=148;
				end
				if(in == 916) begin
					state<=16;
					out<=149;
				end
				if(in == 917) begin
					state<=16;
					out<=150;
				end
				if(in == 918) begin
					state<=16;
					out<=151;
				end
				if(in == 919) begin
					state<=16;
					out<=152;
				end
				if(in == 920) begin
					state<=16;
					out<=153;
				end
				if(in == 921) begin
					state<=16;
					out<=154;
				end
				if(in == 922) begin
					state<=16;
					out<=155;
				end
				if(in == 923) begin
					state<=16;
					out<=156;
				end
				if(in == 924) begin
					state<=16;
					out<=157;
				end
				if(in == 925) begin
					state<=16;
					out<=158;
				end
				if(in == 926) begin
					state<=16;
					out<=159;
				end
				if(in == 927) begin
					state<=16;
					out<=160;
				end
				if(in == 928) begin
					state<=16;
					out<=161;
				end
			end
			2: begin
				if(in == 0) begin
					state<=3;
					out<=162;
				end
				if(in == 1) begin
					state<=1;
					out<=163;
				end
				if(in == 2) begin
					state<=2;
					out<=164;
				end
				if(in == 3) begin
					state<=3;
					out<=165;
				end
				if(in == 4) begin
					state<=2;
					out<=166;
				end
				if(in == 5) begin
					state<=3;
					out<=167;
				end
				if(in == 6) begin
					state<=2;
					out<=168;
				end
				if(in == 7) begin
					state<=2;
					out<=169;
				end
				if(in == 8) begin
					state<=2;
					out<=170;
				end
				if(in == 9) begin
					state<=2;
					out<=171;
				end
				if(in == 10) begin
					state<=2;
					out<=172;
				end
				if(in == 11) begin
					state<=2;
					out<=173;
				end
				if(in == 12) begin
					state<=2;
					out<=174;
				end
				if(in == 13) begin
					state<=2;
					out<=175;
				end
				if(in == 14) begin
					state<=2;
					out<=176;
				end
				if(in == 15) begin
					state<=2;
					out<=177;
				end
				if(in == 16) begin
					state<=2;
					out<=178;
				end
				if(in == 17) begin
					state<=2;
					out<=179;
				end
				if(in == 18) begin
					state<=2;
					out<=180;
				end
				if(in == 19) begin
					state<=2;
					out<=181;
				end
				if(in == 20) begin
					state<=2;
					out<=182;
				end
				if(in == 21) begin
					state<=2;
					out<=183;
				end
				if(in == 22) begin
					state<=2;
					out<=184;
				end
				if(in == 23) begin
					state<=2;
					out<=185;
				end
				if(in == 24) begin
					state<=2;
					out<=186;
				end
				if(in == 25) begin
					state<=2;
					out<=187;
				end
				if(in == 26) begin
					state<=2;
					out<=188;
				end
				if(in == 27) begin
					state<=2;
					out<=189;
				end
				if(in == 28) begin
					state<=2;
					out<=190;
				end
				if(in == 29) begin
					state<=2;
					out<=191;
				end
				if(in == 30) begin
					state<=2;
					out<=192;
				end
				if(in == 31) begin
					state<=2;
					out<=193;
				end
				if(in == 32) begin
					state<=2;
					out<=194;
				end
				if(in == 33) begin
					state<=2;
					out<=195;
				end
				if(in == 34) begin
					state<=2;
					out<=196;
				end
				if(in == 35) begin
					state<=2;
					out<=197;
				end
				if(in == 36) begin
					state<=2;
					out<=198;
				end
				if(in == 37) begin
					state<=2;
					out<=199;
				end
				if(in == 38) begin
					state<=2;
					out<=200;
				end
				if(in == 39) begin
					state<=2;
					out<=201;
				end
				if(in == 40) begin
					state<=2;
					out<=202;
				end
				if(in == 41) begin
					state<=2;
					out<=203;
				end
				if(in == 42) begin
					state<=2;
					out<=204;
				end
				if(in == 43) begin
					state<=2;
					out<=205;
				end
				if(in == 44) begin
					state<=2;
					out<=206;
				end
				if(in == 45) begin
					state<=2;
					out<=207;
				end
				if(in == 46) begin
					state<=2;
					out<=208;
				end
				if(in == 47) begin
					state<=2;
					out<=209;
				end
				if(in == 48) begin
					state<=2;
					out<=210;
				end
				if(in == 49) begin
					state<=2;
					out<=211;
				end
				if(in == 50) begin
					state<=2;
					out<=212;
				end
				if(in == 51) begin
					state<=2;
					out<=213;
				end
				if(in == 52) begin
					state<=2;
					out<=214;
				end
				if(in == 53) begin
					state<=3;
					out<=215;
				end
				if(in == 54) begin
					state<=2;
					out<=216;
				end
				if(in == 55) begin
					state<=3;
					out<=217;
				end
				if(in == 56) begin
					state<=2;
					out<=218;
				end
				if(in == 57) begin
					state<=3;
					out<=219;
				end
				if(in == 58) begin
					state<=2;
					out<=220;
				end
				if(in == 59) begin
					state<=2;
					out<=221;
				end
				if(in == 60) begin
					state<=2;
					out<=222;
				end
				if(in == 61) begin
					state<=2;
					out<=223;
				end
				if(in == 62) begin
					state<=2;
					out<=224;
				end
				if(in == 63) begin
					state<=2;
					out<=225;
				end
				if(in == 64) begin
					state<=2;
					out<=226;
				end
				if(in == 65) begin
					state<=2;
					out<=227;
				end
				if(in == 66) begin
					state<=2;
					out<=228;
				end
				if(in == 67) begin
					state<=2;
					out<=229;
				end
				if(in == 68) begin
					state<=2;
					out<=230;
				end
				if(in == 69) begin
					state<=2;
					out<=231;
				end
				if(in == 70) begin
					state<=2;
					out<=232;
				end
				if(in == 71) begin
					state<=2;
					out<=233;
				end
				if(in == 72) begin
					state<=2;
					out<=234;
				end
				if(in == 73) begin
					state<=2;
					out<=235;
				end
				if(in == 74) begin
					state<=2;
					out<=236;
				end
				if(in == 75) begin
					state<=2;
					out<=237;
				end
				if(in == 76) begin
					state<=2;
					out<=238;
				end
				if(in == 77) begin
					state<=2;
					out<=239;
				end
				if(in == 78) begin
					state<=2;
					out<=240;
				end
				if(in == 79) begin
					state<=2;
					out<=241;
				end
				if(in == 80) begin
					state<=2;
					out<=242;
				end
				if(in == 81) begin
					state<=2;
					out<=243;
				end
				if(in == 82) begin
					state<=2;
					out<=244;
				end
				if(in == 83) begin
					state<=2;
					out<=245;
				end
				if(in == 84) begin
					state<=2;
					out<=246;
				end
				if(in == 85) begin
					state<=2;
					out<=247;
				end
				if(in == 86) begin
					state<=2;
					out<=248;
				end
				if(in == 87) begin
					state<=2;
					out<=249;
				end
				if(in == 88) begin
					state<=2;
					out<=250;
				end
				if(in == 89) begin
					state<=2;
					out<=251;
				end
				if(in == 90) begin
					state<=2;
					out<=252;
				end
				if(in == 91) begin
					state<=2;
					out<=253;
				end
				if(in == 92) begin
					state<=2;
					out<=254;
				end
				if(in == 93) begin
					state<=2;
					out<=255;
				end
				if(in == 94) begin
					state<=2;
					out<=0;
				end
				if(in == 95) begin
					state<=2;
					out<=1;
				end
				if(in == 96) begin
					state<=2;
					out<=2;
				end
				if(in == 97) begin
					state<=2;
					out<=3;
				end
				if(in == 98) begin
					state<=2;
					out<=4;
				end
				if(in == 99) begin
					state<=2;
					out<=5;
				end
				if(in == 100) begin
					state<=2;
					out<=6;
				end
				if(in == 101) begin
					state<=2;
					out<=7;
				end
				if(in == 102) begin
					state<=2;
					out<=8;
				end
				if(in == 103) begin
					state<=2;
					out<=9;
				end
				if(in == 104) begin
					state<=2;
					out<=10;
				end
				if(in == 105) begin
					state<=3;
					out<=11;
				end
				if(in == 106) begin
					state<=2;
					out<=12;
				end
				if(in == 107) begin
					state<=3;
					out<=13;
				end
				if(in == 108) begin
					state<=2;
					out<=14;
				end
				if(in == 109) begin
					state<=3;
					out<=15;
				end
				if(in == 110) begin
					state<=2;
					out<=16;
				end
				if(in == 111) begin
					state<=3;
					out<=17;
				end
				if(in == 112) begin
					state<=2;
					out<=18;
				end
				if(in == 113) begin
					state<=3;
					out<=19;
				end
				if(in == 114) begin
					state<=2;
					out<=20;
				end
				if(in == 115) begin
					state<=3;
					out<=21;
				end
				if(in == 116) begin
					state<=2;
					out<=22;
				end
				if(in == 117) begin
					state<=3;
					out<=23;
				end
				if(in == 118) begin
					state<=2;
					out<=24;
				end
				if(in == 119) begin
					state<=3;
					out<=25;
				end
				if(in == 120) begin
					state<=2;
					out<=26;
				end
				if(in == 121) begin
					state<=3;
					out<=27;
				end
				if(in == 122) begin
					state<=2;
					out<=28;
				end
				if(in == 123) begin
					state<=2;
					out<=29;
				end
				if(in == 124) begin
					state<=2;
					out<=30;
				end
				if(in == 125) begin
					state<=2;
					out<=31;
				end
				if(in == 126) begin
					state<=2;
					out<=32;
				end
				if(in == 127) begin
					state<=2;
					out<=33;
				end
				if(in == 128) begin
					state<=2;
					out<=34;
				end
				if(in == 129) begin
					state<=2;
					out<=35;
				end
				if(in == 130) begin
					state<=2;
					out<=36;
				end
				if(in == 131) begin
					state<=2;
					out<=37;
				end
				if(in == 132) begin
					state<=2;
					out<=38;
				end
				if(in == 133) begin
					state<=2;
					out<=39;
				end
				if(in == 134) begin
					state<=2;
					out<=40;
				end
				if(in == 135) begin
					state<=2;
					out<=41;
				end
				if(in == 136) begin
					state<=2;
					out<=42;
				end
				if(in == 137) begin
					state<=2;
					out<=43;
				end
				if(in == 138) begin
					state<=2;
					out<=44;
				end
				if(in == 139) begin
					state<=2;
					out<=45;
				end
				if(in == 140) begin
					state<=2;
					out<=46;
				end
				if(in == 141) begin
					state<=2;
					out<=47;
				end
				if(in == 142) begin
					state<=2;
					out<=48;
				end
				if(in == 143) begin
					state<=2;
					out<=49;
				end
				if(in == 144) begin
					state<=2;
					out<=50;
				end
				if(in == 145) begin
					state<=2;
					out<=51;
				end
				if(in == 146) begin
					state<=2;
					out<=52;
				end
				if(in == 147) begin
					state<=2;
					out<=53;
				end
				if(in == 148) begin
					state<=2;
					out<=54;
				end
				if(in == 149) begin
					state<=2;
					out<=55;
				end
				if(in == 150) begin
					state<=2;
					out<=56;
				end
				if(in == 151) begin
					state<=2;
					out<=57;
				end
				if(in == 152) begin
					state<=2;
					out<=58;
				end
				if(in == 153) begin
					state<=2;
					out<=59;
				end
				if(in == 154) begin
					state<=2;
					out<=60;
				end
				if(in == 155) begin
					state<=2;
					out<=61;
				end
				if(in == 156) begin
					state<=2;
					out<=62;
				end
				if(in == 157) begin
					state<=2;
					out<=63;
				end
				if(in == 158) begin
					state<=2;
					out<=64;
				end
				if(in == 159) begin
					state<=2;
					out<=65;
				end
				if(in == 160) begin
					state<=2;
					out<=66;
				end
				if(in == 161) begin
					state<=2;
					out<=67;
				end
				if(in == 162) begin
					state<=2;
					out<=68;
				end
				if(in == 163) begin
					state<=2;
					out<=69;
				end
				if(in == 164) begin
					state<=2;
					out<=70;
				end
				if(in == 165) begin
					state<=2;
					out<=71;
				end
				if(in == 166) begin
					state<=2;
					out<=72;
				end
				if(in == 167) begin
					state<=2;
					out<=73;
				end
				if(in == 168) begin
					state<=2;
					out<=74;
				end
				if(in == 169) begin
					state<=3;
					out<=75;
				end
				if(in == 170) begin
					state<=2;
					out<=76;
				end
				if(in == 171) begin
					state<=3;
					out<=77;
				end
				if(in == 172) begin
					state<=2;
					out<=78;
				end
				if(in == 173) begin
					state<=3;
					out<=79;
				end
				if(in == 174) begin
					state<=2;
					out<=80;
				end
				if(in == 175) begin
					state<=2;
					out<=81;
				end
				if(in == 176) begin
					state<=2;
					out<=82;
				end
				if(in == 177) begin
					state<=2;
					out<=83;
				end
				if(in == 178) begin
					state<=2;
					out<=84;
				end
				if(in == 179) begin
					state<=2;
					out<=85;
				end
				if(in == 180) begin
					state<=2;
					out<=86;
				end
				if(in == 181) begin
					state<=2;
					out<=87;
				end
				if(in == 182) begin
					state<=2;
					out<=88;
				end
				if(in == 183) begin
					state<=2;
					out<=89;
				end
				if(in == 184) begin
					state<=2;
					out<=90;
				end
				if(in == 185) begin
					state<=2;
					out<=91;
				end
				if(in == 186) begin
					state<=2;
					out<=92;
				end
				if(in == 187) begin
					state<=2;
					out<=93;
				end
				if(in == 188) begin
					state<=2;
					out<=94;
				end
				if(in == 189) begin
					state<=2;
					out<=95;
				end
				if(in == 190) begin
					state<=2;
					out<=96;
				end
				if(in == 191) begin
					state<=2;
					out<=97;
				end
				if(in == 192) begin
					state<=2;
					out<=98;
				end
				if(in == 193) begin
					state<=2;
					out<=99;
				end
				if(in == 194) begin
					state<=2;
					out<=100;
				end
				if(in == 195) begin
					state<=2;
					out<=101;
				end
				if(in == 196) begin
					state<=2;
					out<=102;
				end
				if(in == 197) begin
					state<=2;
					out<=103;
				end
				if(in == 198) begin
					state<=2;
					out<=104;
				end
				if(in == 199) begin
					state<=2;
					out<=105;
				end
				if(in == 200) begin
					state<=2;
					out<=106;
				end
				if(in == 201) begin
					state<=2;
					out<=107;
				end
				if(in == 202) begin
					state<=2;
					out<=108;
				end
				if(in == 203) begin
					state<=2;
					out<=109;
				end
				if(in == 204) begin
					state<=2;
					out<=110;
				end
				if(in == 205) begin
					state<=2;
					out<=111;
				end
				if(in == 206) begin
					state<=2;
					out<=112;
				end
				if(in == 207) begin
					state<=2;
					out<=113;
				end
				if(in == 208) begin
					state<=2;
					out<=114;
				end
				if(in == 209) begin
					state<=2;
					out<=115;
				end
				if(in == 210) begin
					state<=2;
					out<=116;
				end
				if(in == 211) begin
					state<=2;
					out<=117;
				end
				if(in == 212) begin
					state<=2;
					out<=118;
				end
				if(in == 213) begin
					state<=2;
					out<=119;
				end
				if(in == 214) begin
					state<=2;
					out<=120;
				end
				if(in == 215) begin
					state<=2;
					out<=121;
				end
				if(in == 216) begin
					state<=2;
					out<=122;
				end
				if(in == 217) begin
					state<=2;
					out<=123;
				end
				if(in == 218) begin
					state<=2;
					out<=124;
				end
				if(in == 219) begin
					state<=2;
					out<=125;
				end
				if(in == 220) begin
					state<=2;
					out<=126;
				end
				if(in == 221) begin
					state<=3;
					out<=127;
				end
				if(in == 222) begin
					state<=2;
					out<=128;
				end
				if(in == 223) begin
					state<=3;
					out<=129;
				end
				if(in == 224) begin
					state<=2;
					out<=130;
				end
				if(in == 225) begin
					state<=3;
					out<=131;
				end
				if(in == 226) begin
					state<=2;
					out<=132;
				end
				if(in == 227) begin
					state<=3;
					out<=133;
				end
				if(in == 228) begin
					state<=2;
					out<=134;
				end
				if(in == 229) begin
					state<=3;
					out<=135;
				end
				if(in == 230) begin
					state<=2;
					out<=136;
				end
				if(in == 231) begin
					state<=3;
					out<=137;
				end
				if(in == 232) begin
					state<=2;
					out<=138;
				end
				if(in == 233) begin
					state<=3;
					out<=139;
				end
				if(in == 234) begin
					state<=2;
					out<=140;
				end
				if(in == 235) begin
					state<=3;
					out<=141;
				end
				if(in == 236) begin
					state<=2;
					out<=142;
				end
				if(in == 237) begin
					state<=3;
					out<=143;
				end
				if(in == 238) begin
					state<=2;
					out<=144;
				end
				if(in == 239) begin
					state<=2;
					out<=145;
				end
				if(in == 240) begin
					state<=2;
					out<=146;
				end
				if(in == 241) begin
					state<=2;
					out<=147;
				end
				if(in == 242) begin
					state<=2;
					out<=148;
				end
				if(in == 243) begin
					state<=2;
					out<=149;
				end
				if(in == 244) begin
					state<=2;
					out<=150;
				end
				if(in == 245) begin
					state<=2;
					out<=151;
				end
				if(in == 246) begin
					state<=2;
					out<=152;
				end
				if(in == 247) begin
					state<=2;
					out<=153;
				end
				if(in == 248) begin
					state<=2;
					out<=154;
				end
				if(in == 249) begin
					state<=2;
					out<=155;
				end
				if(in == 250) begin
					state<=2;
					out<=156;
				end
				if(in == 251) begin
					state<=2;
					out<=157;
				end
				if(in == 252) begin
					state<=2;
					out<=158;
				end
				if(in == 253) begin
					state<=2;
					out<=159;
				end
				if(in == 254) begin
					state<=2;
					out<=160;
				end
				if(in == 255) begin
					state<=2;
					out<=161;
				end
				if(in == 256) begin
					state<=2;
					out<=162;
				end
				if(in == 257) begin
					state<=2;
					out<=163;
				end
				if(in == 258) begin
					state<=2;
					out<=164;
				end
				if(in == 259) begin
					state<=2;
					out<=165;
				end
				if(in == 260) begin
					state<=2;
					out<=166;
				end
				if(in == 261) begin
					state<=2;
					out<=167;
				end
				if(in == 262) begin
					state<=2;
					out<=168;
				end
				if(in == 263) begin
					state<=2;
					out<=169;
				end
				if(in == 264) begin
					state<=2;
					out<=170;
				end
				if(in == 265) begin
					state<=2;
					out<=171;
				end
				if(in == 266) begin
					state<=2;
					out<=172;
				end
				if(in == 267) begin
					state<=2;
					out<=173;
				end
				if(in == 268) begin
					state<=2;
					out<=174;
				end
				if(in == 269) begin
					state<=2;
					out<=175;
				end
				if(in == 270) begin
					state<=2;
					out<=176;
				end
				if(in == 271) begin
					state<=2;
					out<=177;
				end
				if(in == 272) begin
					state<=2;
					out<=178;
				end
				if(in == 273) begin
					state<=2;
					out<=179;
				end
				if(in == 274) begin
					state<=2;
					out<=180;
				end
				if(in == 275) begin
					state<=2;
					out<=181;
				end
				if(in == 276) begin
					state<=2;
					out<=182;
				end
				if(in == 277) begin
					state<=2;
					out<=183;
				end
				if(in == 278) begin
					state<=2;
					out<=184;
				end
				if(in == 279) begin
					state<=2;
					out<=185;
				end
				if(in == 280) begin
					state<=2;
					out<=186;
				end
				if(in == 281) begin
					state<=2;
					out<=187;
				end
				if(in == 282) begin
					state<=2;
					out<=188;
				end
				if(in == 283) begin
					state<=2;
					out<=189;
				end
				if(in == 284) begin
					state<=2;
					out<=190;
				end
				if(in == 285) begin
					state<=3;
					out<=191;
				end
				if(in == 286) begin
					state<=2;
					out<=192;
				end
				if(in == 287) begin
					state<=3;
					out<=193;
				end
				if(in == 288) begin
					state<=2;
					out<=194;
				end
				if(in == 289) begin
					state<=3;
					out<=195;
				end
				if(in == 290) begin
					state<=2;
					out<=196;
				end
				if(in == 291) begin
					state<=2;
					out<=197;
				end
				if(in == 292) begin
					state<=2;
					out<=198;
				end
				if(in == 293) begin
					state<=2;
					out<=199;
				end
				if(in == 294) begin
					state<=2;
					out<=200;
				end
				if(in == 295) begin
					state<=2;
					out<=201;
				end
				if(in == 296) begin
					state<=2;
					out<=202;
				end
				if(in == 297) begin
					state<=2;
					out<=203;
				end
				if(in == 298) begin
					state<=2;
					out<=204;
				end
				if(in == 299) begin
					state<=2;
					out<=205;
				end
				if(in == 300) begin
					state<=2;
					out<=206;
				end
				if(in == 301) begin
					state<=2;
					out<=207;
				end
				if(in == 302) begin
					state<=2;
					out<=208;
				end
				if(in == 303) begin
					state<=2;
					out<=209;
				end
				if(in == 304) begin
					state<=2;
					out<=210;
				end
				if(in == 305) begin
					state<=2;
					out<=211;
				end
				if(in == 306) begin
					state<=2;
					out<=212;
				end
				if(in == 307) begin
					state<=2;
					out<=213;
				end
				if(in == 308) begin
					state<=2;
					out<=214;
				end
				if(in == 309) begin
					state<=2;
					out<=215;
				end
				if(in == 310) begin
					state<=2;
					out<=216;
				end
				if(in == 311) begin
					state<=2;
					out<=217;
				end
				if(in == 312) begin
					state<=2;
					out<=218;
				end
				if(in == 313) begin
					state<=2;
					out<=219;
				end
				if(in == 314) begin
					state<=2;
					out<=220;
				end
				if(in == 315) begin
					state<=2;
					out<=221;
				end
				if(in == 316) begin
					state<=2;
					out<=222;
				end
				if(in == 317) begin
					state<=2;
					out<=223;
				end
				if(in == 318) begin
					state<=2;
					out<=224;
				end
				if(in == 319) begin
					state<=2;
					out<=225;
				end
				if(in == 320) begin
					state<=2;
					out<=226;
				end
				if(in == 321) begin
					state<=2;
					out<=227;
				end
				if(in == 322) begin
					state<=2;
					out<=228;
				end
				if(in == 323) begin
					state<=2;
					out<=229;
				end
				if(in == 324) begin
					state<=2;
					out<=230;
				end
				if(in == 325) begin
					state<=2;
					out<=231;
				end
				if(in == 326) begin
					state<=2;
					out<=232;
				end
				if(in == 327) begin
					state<=2;
					out<=233;
				end
				if(in == 328) begin
					state<=2;
					out<=234;
				end
				if(in == 329) begin
					state<=2;
					out<=235;
				end
				if(in == 330) begin
					state<=2;
					out<=236;
				end
				if(in == 331) begin
					state<=2;
					out<=237;
				end
				if(in == 332) begin
					state<=2;
					out<=238;
				end
				if(in == 333) begin
					state<=2;
					out<=239;
				end
				if(in == 334) begin
					state<=2;
					out<=240;
				end
				if(in == 335) begin
					state<=2;
					out<=241;
				end
				if(in == 336) begin
					state<=2;
					out<=242;
				end
				if(in == 337) begin
					state<=3;
					out<=243;
				end
				if(in == 338) begin
					state<=2;
					out<=244;
				end
				if(in == 339) begin
					state<=3;
					out<=245;
				end
				if(in == 340) begin
					state<=2;
					out<=246;
				end
				if(in == 341) begin
					state<=3;
					out<=247;
				end
				if(in == 342) begin
					state<=2;
					out<=248;
				end
				if(in == 343) begin
					state<=3;
					out<=249;
				end
				if(in == 344) begin
					state<=2;
					out<=250;
				end
				if(in == 345) begin
					state<=3;
					out<=251;
				end
				if(in == 346) begin
					state<=2;
					out<=252;
				end
				if(in == 347) begin
					state<=3;
					out<=253;
				end
				if(in == 348) begin
					state<=2;
					out<=254;
				end
				if(in == 349) begin
					state<=3;
					out<=255;
				end
				if(in == 350) begin
					state<=2;
					out<=0;
				end
				if(in == 351) begin
					state<=3;
					out<=1;
				end
				if(in == 352) begin
					state<=2;
					out<=2;
				end
				if(in == 353) begin
					state<=3;
					out<=3;
				end
				if(in == 354) begin
					state<=2;
					out<=4;
				end
				if(in == 355) begin
					state<=2;
					out<=5;
				end
				if(in == 356) begin
					state<=2;
					out<=6;
				end
				if(in == 357) begin
					state<=2;
					out<=7;
				end
				if(in == 358) begin
					state<=2;
					out<=8;
				end
				if(in == 359) begin
					state<=2;
					out<=9;
				end
				if(in == 360) begin
					state<=2;
					out<=10;
				end
				if(in == 361) begin
					state<=2;
					out<=11;
				end
				if(in == 362) begin
					state<=2;
					out<=12;
				end
				if(in == 363) begin
					state<=2;
					out<=13;
				end
				if(in == 364) begin
					state<=2;
					out<=14;
				end
				if(in == 365) begin
					state<=2;
					out<=15;
				end
				if(in == 366) begin
					state<=2;
					out<=16;
				end
				if(in == 367) begin
					state<=2;
					out<=17;
				end
				if(in == 368) begin
					state<=2;
					out<=18;
				end
				if(in == 369) begin
					state<=2;
					out<=19;
				end
				if(in == 370) begin
					state<=2;
					out<=20;
				end
				if(in == 371) begin
					state<=2;
					out<=21;
				end
				if(in == 372) begin
					state<=2;
					out<=22;
				end
				if(in == 373) begin
					state<=2;
					out<=23;
				end
				if(in == 374) begin
					state<=2;
					out<=24;
				end
				if(in == 375) begin
					state<=2;
					out<=25;
				end
				if(in == 376) begin
					state<=2;
					out<=26;
				end
				if(in == 377) begin
					state<=2;
					out<=27;
				end
				if(in == 378) begin
					state<=2;
					out<=28;
				end
				if(in == 379) begin
					state<=2;
					out<=29;
				end
				if(in == 380) begin
					state<=2;
					out<=30;
				end
				if(in == 381) begin
					state<=2;
					out<=31;
				end
				if(in == 382) begin
					state<=2;
					out<=32;
				end
				if(in == 383) begin
					state<=2;
					out<=33;
				end
				if(in == 384) begin
					state<=2;
					out<=34;
				end
				if(in == 385) begin
					state<=2;
					out<=35;
				end
				if(in == 386) begin
					state<=2;
					out<=36;
				end
				if(in == 387) begin
					state<=2;
					out<=37;
				end
				if(in == 388) begin
					state<=2;
					out<=38;
				end
				if(in == 389) begin
					state<=2;
					out<=39;
				end
				if(in == 390) begin
					state<=2;
					out<=40;
				end
				if(in == 391) begin
					state<=2;
					out<=41;
				end
				if(in == 392) begin
					state<=2;
					out<=42;
				end
				if(in == 393) begin
					state<=2;
					out<=43;
				end
				if(in == 394) begin
					state<=2;
					out<=44;
				end
				if(in == 395) begin
					state<=2;
					out<=45;
				end
				if(in == 396) begin
					state<=2;
					out<=46;
				end
				if(in == 397) begin
					state<=2;
					out<=47;
				end
				if(in == 398) begin
					state<=2;
					out<=48;
				end
				if(in == 399) begin
					state<=2;
					out<=49;
				end
				if(in == 400) begin
					state<=2;
					out<=50;
				end
				if(in == 401) begin
					state<=3;
					out<=51;
				end
				if(in == 402) begin
					state<=2;
					out<=52;
				end
				if(in == 403) begin
					state<=3;
					out<=53;
				end
				if(in == 404) begin
					state<=2;
					out<=54;
				end
				if(in == 405) begin
					state<=3;
					out<=55;
				end
				if(in == 406) begin
					state<=2;
					out<=56;
				end
				if(in == 407) begin
					state<=2;
					out<=57;
				end
				if(in == 408) begin
					state<=2;
					out<=58;
				end
				if(in == 409) begin
					state<=2;
					out<=59;
				end
				if(in == 410) begin
					state<=2;
					out<=60;
				end
				if(in == 411) begin
					state<=2;
					out<=61;
				end
				if(in == 412) begin
					state<=2;
					out<=62;
				end
				if(in == 413) begin
					state<=2;
					out<=63;
				end
				if(in == 414) begin
					state<=2;
					out<=64;
				end
				if(in == 415) begin
					state<=2;
					out<=65;
				end
				if(in == 416) begin
					state<=2;
					out<=66;
				end
				if(in == 417) begin
					state<=2;
					out<=67;
				end
				if(in == 418) begin
					state<=2;
					out<=68;
				end
				if(in == 419) begin
					state<=2;
					out<=69;
				end
				if(in == 420) begin
					state<=2;
					out<=70;
				end
				if(in == 421) begin
					state<=2;
					out<=71;
				end
				if(in == 422) begin
					state<=2;
					out<=72;
				end
				if(in == 423) begin
					state<=2;
					out<=73;
				end
				if(in == 424) begin
					state<=2;
					out<=74;
				end
				if(in == 425) begin
					state<=2;
					out<=75;
				end
				if(in == 426) begin
					state<=2;
					out<=76;
				end
				if(in == 427) begin
					state<=2;
					out<=77;
				end
				if(in == 428) begin
					state<=2;
					out<=78;
				end
				if(in == 429) begin
					state<=2;
					out<=79;
				end
				if(in == 430) begin
					state<=2;
					out<=80;
				end
				if(in == 431) begin
					state<=2;
					out<=81;
				end
				if(in == 432) begin
					state<=2;
					out<=82;
				end
				if(in == 433) begin
					state<=2;
					out<=83;
				end
				if(in == 434) begin
					state<=2;
					out<=84;
				end
				if(in == 435) begin
					state<=2;
					out<=85;
				end
				if(in == 436) begin
					state<=2;
					out<=86;
				end
				if(in == 437) begin
					state<=2;
					out<=87;
				end
				if(in == 438) begin
					state<=2;
					out<=88;
				end
				if(in == 439) begin
					state<=2;
					out<=89;
				end
				if(in == 440) begin
					state<=2;
					out<=90;
				end
				if(in == 441) begin
					state<=2;
					out<=91;
				end
				if(in == 442) begin
					state<=2;
					out<=92;
				end
				if(in == 443) begin
					state<=2;
					out<=93;
				end
				if(in == 444) begin
					state<=2;
					out<=94;
				end
				if(in == 445) begin
					state<=2;
					out<=95;
				end
				if(in == 446) begin
					state<=2;
					out<=96;
				end
				if(in == 447) begin
					state<=2;
					out<=97;
				end
				if(in == 448) begin
					state<=2;
					out<=98;
				end
				if(in == 449) begin
					state<=2;
					out<=99;
				end
				if(in == 450) begin
					state<=2;
					out<=100;
				end
				if(in == 451) begin
					state<=2;
					out<=101;
				end
				if(in == 452) begin
					state<=2;
					out<=102;
				end
				if(in == 453) begin
					state<=3;
					out<=103;
				end
				if(in == 454) begin
					state<=2;
					out<=104;
				end
				if(in == 455) begin
					state<=3;
					out<=105;
				end
				if(in == 456) begin
					state<=2;
					out<=106;
				end
				if(in == 457) begin
					state<=3;
					out<=107;
				end
				if(in == 458) begin
					state<=2;
					out<=108;
				end
				if(in == 459) begin
					state<=3;
					out<=109;
				end
				if(in == 460) begin
					state<=2;
					out<=110;
				end
				if(in == 461) begin
					state<=3;
					out<=111;
				end
				if(in == 462) begin
					state<=2;
					out<=112;
				end
				if(in == 463) begin
					state<=3;
					out<=113;
				end
				if(in == 464) begin
					state<=2;
					out<=114;
				end
				if(in == 465) begin
					state<=3;
					out<=115;
				end
				if(in == 466) begin
					state<=2;
					out<=116;
				end
				if(in == 467) begin
					state<=3;
					out<=117;
				end
				if(in == 468) begin
					state<=2;
					out<=118;
				end
				if(in == 469) begin
					state<=3;
					out<=119;
				end
				if(in == 470) begin
					state<=2;
					out<=120;
				end
				if(in == 471) begin
					state<=2;
					out<=121;
				end
				if(in == 472) begin
					state<=2;
					out<=122;
				end
				if(in == 473) begin
					state<=2;
					out<=123;
				end
				if(in == 474) begin
					state<=2;
					out<=124;
				end
				if(in == 475) begin
					state<=2;
					out<=125;
				end
				if(in == 476) begin
					state<=2;
					out<=126;
				end
				if(in == 477) begin
					state<=2;
					out<=127;
				end
				if(in == 478) begin
					state<=2;
					out<=128;
				end
				if(in == 479) begin
					state<=2;
					out<=129;
				end
				if(in == 480) begin
					state<=2;
					out<=130;
				end
				if(in == 481) begin
					state<=2;
					out<=131;
				end
				if(in == 482) begin
					state<=2;
					out<=132;
				end
				if(in == 483) begin
					state<=2;
					out<=133;
				end
				if(in == 484) begin
					state<=2;
					out<=134;
				end
				if(in == 485) begin
					state<=2;
					out<=135;
				end
				if(in == 486) begin
					state<=2;
					out<=136;
				end
				if(in == 487) begin
					state<=2;
					out<=137;
				end
				if(in == 488) begin
					state<=2;
					out<=138;
				end
				if(in == 489) begin
					state<=2;
					out<=139;
				end
				if(in == 490) begin
					state<=2;
					out<=140;
				end
				if(in == 491) begin
					state<=2;
					out<=141;
				end
				if(in == 492) begin
					state<=2;
					out<=142;
				end
				if(in == 493) begin
					state<=2;
					out<=143;
				end
				if(in == 494) begin
					state<=2;
					out<=144;
				end
				if(in == 495) begin
					state<=2;
					out<=145;
				end
				if(in == 496) begin
					state<=2;
					out<=146;
				end
				if(in == 497) begin
					state<=2;
					out<=147;
				end
				if(in == 498) begin
					state<=2;
					out<=148;
				end
				if(in == 499) begin
					state<=2;
					out<=149;
				end
				if(in == 500) begin
					state<=2;
					out<=150;
				end
				if(in == 501) begin
					state<=2;
					out<=151;
				end
				if(in == 502) begin
					state<=2;
					out<=152;
				end
				if(in == 503) begin
					state<=2;
					out<=153;
				end
				if(in == 504) begin
					state<=2;
					out<=154;
				end
				if(in == 505) begin
					state<=2;
					out<=155;
				end
				if(in == 506) begin
					state<=2;
					out<=156;
				end
				if(in == 507) begin
					state<=2;
					out<=157;
				end
				if(in == 508) begin
					state<=2;
					out<=158;
				end
				if(in == 509) begin
					state<=2;
					out<=159;
				end
				if(in == 510) begin
					state<=2;
					out<=160;
				end
				if(in == 511) begin
					state<=2;
					out<=161;
				end
				if(in == 512) begin
					state<=2;
					out<=162;
				end
				if(in == 513) begin
					state<=2;
					out<=163;
				end
				if(in == 514) begin
					state<=2;
					out<=164;
				end
				if(in == 515) begin
					state<=2;
					out<=165;
				end
				if(in == 516) begin
					state<=2;
					out<=166;
				end
				if(in == 517) begin
					state<=3;
					out<=167;
				end
				if(in == 518) begin
					state<=2;
					out<=168;
				end
				if(in == 519) begin
					state<=3;
					out<=169;
				end
				if(in == 520) begin
					state<=2;
					out<=170;
				end
				if(in == 521) begin
					state<=3;
					out<=171;
				end
				if(in == 522) begin
					state<=2;
					out<=172;
				end
				if(in == 523) begin
					state<=2;
					out<=173;
				end
				if(in == 524) begin
					state<=2;
					out<=174;
				end
				if(in == 525) begin
					state<=2;
					out<=175;
				end
				if(in == 526) begin
					state<=2;
					out<=176;
				end
				if(in == 527) begin
					state<=2;
					out<=177;
				end
				if(in == 528) begin
					state<=2;
					out<=178;
				end
				if(in == 529) begin
					state<=2;
					out<=179;
				end
				if(in == 530) begin
					state<=2;
					out<=180;
				end
				if(in == 531) begin
					state<=2;
					out<=181;
				end
				if(in == 532) begin
					state<=2;
					out<=182;
				end
				if(in == 533) begin
					state<=2;
					out<=183;
				end
				if(in == 534) begin
					state<=2;
					out<=184;
				end
				if(in == 535) begin
					state<=2;
					out<=185;
				end
				if(in == 536) begin
					state<=2;
					out<=186;
				end
				if(in == 537) begin
					state<=2;
					out<=187;
				end
				if(in == 538) begin
					state<=2;
					out<=188;
				end
				if(in == 539) begin
					state<=2;
					out<=189;
				end
				if(in == 540) begin
					state<=2;
					out<=190;
				end
				if(in == 541) begin
					state<=2;
					out<=191;
				end
				if(in == 542) begin
					state<=2;
					out<=192;
				end
				if(in == 543) begin
					state<=2;
					out<=193;
				end
				if(in == 544) begin
					state<=2;
					out<=194;
				end
				if(in == 545) begin
					state<=2;
					out<=195;
				end
				if(in == 546) begin
					state<=2;
					out<=196;
				end
				if(in == 547) begin
					state<=2;
					out<=197;
				end
				if(in == 548) begin
					state<=2;
					out<=198;
				end
				if(in == 549) begin
					state<=2;
					out<=199;
				end
				if(in == 550) begin
					state<=2;
					out<=200;
				end
				if(in == 551) begin
					state<=2;
					out<=201;
				end
				if(in == 552) begin
					state<=2;
					out<=202;
				end
				if(in == 553) begin
					state<=2;
					out<=203;
				end
				if(in == 554) begin
					state<=2;
					out<=204;
				end
				if(in == 555) begin
					state<=2;
					out<=205;
				end
				if(in == 556) begin
					state<=2;
					out<=206;
				end
				if(in == 557) begin
					state<=2;
					out<=207;
				end
				if(in == 558) begin
					state<=2;
					out<=208;
				end
				if(in == 559) begin
					state<=2;
					out<=209;
				end
				if(in == 560) begin
					state<=2;
					out<=210;
				end
				if(in == 561) begin
					state<=2;
					out<=211;
				end
				if(in == 562) begin
					state<=2;
					out<=212;
				end
				if(in == 563) begin
					state<=2;
					out<=213;
				end
				if(in == 564) begin
					state<=2;
					out<=214;
				end
				if(in == 565) begin
					state<=2;
					out<=215;
				end
				if(in == 566) begin
					state<=2;
					out<=216;
				end
				if(in == 567) begin
					state<=2;
					out<=217;
				end
				if(in == 568) begin
					state<=2;
					out<=218;
				end
				if(in == 569) begin
					state<=3;
					out<=219;
				end
				if(in == 570) begin
					state<=2;
					out<=220;
				end
				if(in == 571) begin
					state<=3;
					out<=221;
				end
				if(in == 572) begin
					state<=2;
					out<=222;
				end
				if(in == 573) begin
					state<=3;
					out<=223;
				end
				if(in == 574) begin
					state<=2;
					out<=224;
				end
				if(in == 575) begin
					state<=3;
					out<=225;
				end
				if(in == 576) begin
					state<=2;
					out<=226;
				end
				if(in == 577) begin
					state<=3;
					out<=227;
				end
				if(in == 578) begin
					state<=2;
					out<=228;
				end
				if(in == 579) begin
					state<=3;
					out<=229;
				end
				if(in == 580) begin
					state<=2;
					out<=230;
				end
				if(in == 581) begin
					state<=3;
					out<=231;
				end
				if(in == 582) begin
					state<=2;
					out<=232;
				end
				if(in == 583) begin
					state<=3;
					out<=233;
				end
				if(in == 584) begin
					state<=2;
					out<=234;
				end
				if(in == 585) begin
					state<=3;
					out<=235;
				end
				if(in == 586) begin
					state<=2;
					out<=236;
				end
				if(in == 587) begin
					state<=2;
					out<=237;
				end
				if(in == 588) begin
					state<=2;
					out<=238;
				end
				if(in == 589) begin
					state<=2;
					out<=239;
				end
				if(in == 590) begin
					state<=2;
					out<=240;
				end
				if(in == 591) begin
					state<=2;
					out<=241;
				end
				if(in == 592) begin
					state<=2;
					out<=242;
				end
				if(in == 593) begin
					state<=2;
					out<=243;
				end
				if(in == 594) begin
					state<=2;
					out<=244;
				end
				if(in == 595) begin
					state<=2;
					out<=245;
				end
				if(in == 596) begin
					state<=2;
					out<=246;
				end
				if(in == 597) begin
					state<=2;
					out<=247;
				end
				if(in == 598) begin
					state<=2;
					out<=248;
				end
				if(in == 599) begin
					state<=2;
					out<=249;
				end
				if(in == 600) begin
					state<=2;
					out<=250;
				end
				if(in == 601) begin
					state<=2;
					out<=251;
				end
				if(in == 602) begin
					state<=2;
					out<=252;
				end
				if(in == 603) begin
					state<=2;
					out<=253;
				end
				if(in == 604) begin
					state<=2;
					out<=254;
				end
				if(in == 605) begin
					state<=2;
					out<=255;
				end
				if(in == 606) begin
					state<=2;
					out<=0;
				end
				if(in == 607) begin
					state<=2;
					out<=1;
				end
				if(in == 608) begin
					state<=2;
					out<=2;
				end
				if(in == 609) begin
					state<=2;
					out<=3;
				end
				if(in == 610) begin
					state<=2;
					out<=4;
				end
				if(in == 611) begin
					state<=2;
					out<=5;
				end
				if(in == 612) begin
					state<=2;
					out<=6;
				end
				if(in == 613) begin
					state<=2;
					out<=7;
				end
				if(in == 614) begin
					state<=2;
					out<=8;
				end
				if(in == 615) begin
					state<=2;
					out<=9;
				end
				if(in == 616) begin
					state<=2;
					out<=10;
				end
				if(in == 617) begin
					state<=2;
					out<=11;
				end
				if(in == 618) begin
					state<=2;
					out<=12;
				end
				if(in == 619) begin
					state<=2;
					out<=13;
				end
				if(in == 620) begin
					state<=2;
					out<=14;
				end
				if(in == 621) begin
					state<=2;
					out<=15;
				end
				if(in == 622) begin
					state<=2;
					out<=16;
				end
				if(in == 623) begin
					state<=2;
					out<=17;
				end
				if(in == 624) begin
					state<=2;
					out<=18;
				end
				if(in == 625) begin
					state<=2;
					out<=19;
				end
				if(in == 626) begin
					state<=2;
					out<=20;
				end
				if(in == 627) begin
					state<=2;
					out<=21;
				end
				if(in == 628) begin
					state<=2;
					out<=22;
				end
				if(in == 629) begin
					state<=2;
					out<=23;
				end
				if(in == 630) begin
					state<=2;
					out<=24;
				end
				if(in == 631) begin
					state<=2;
					out<=25;
				end
				if(in == 632) begin
					state<=2;
					out<=26;
				end
				if(in == 633) begin
					state<=3;
					out<=27;
				end
				if(in == 634) begin
					state<=2;
					out<=28;
				end
				if(in == 635) begin
					state<=3;
					out<=29;
				end
				if(in == 636) begin
					state<=2;
					out<=30;
				end
				if(in == 637) begin
					state<=3;
					out<=31;
				end
				if(in == 638) begin
					state<=2;
					out<=32;
				end
				if(in == 639) begin
					state<=2;
					out<=33;
				end
				if(in == 640) begin
					state<=2;
					out<=34;
				end
				if(in == 641) begin
					state<=2;
					out<=35;
				end
				if(in == 642) begin
					state<=2;
					out<=36;
				end
				if(in == 643) begin
					state<=2;
					out<=37;
				end
				if(in == 644) begin
					state<=2;
					out<=38;
				end
				if(in == 645) begin
					state<=2;
					out<=39;
				end
				if(in == 646) begin
					state<=2;
					out<=40;
				end
				if(in == 647) begin
					state<=2;
					out<=41;
				end
				if(in == 648) begin
					state<=2;
					out<=42;
				end
				if(in == 649) begin
					state<=2;
					out<=43;
				end
				if(in == 650) begin
					state<=2;
					out<=44;
				end
				if(in == 651) begin
					state<=2;
					out<=45;
				end
				if(in == 652) begin
					state<=2;
					out<=46;
				end
				if(in == 653) begin
					state<=2;
					out<=47;
				end
				if(in == 654) begin
					state<=2;
					out<=48;
				end
				if(in == 655) begin
					state<=2;
					out<=49;
				end
				if(in == 656) begin
					state<=2;
					out<=50;
				end
				if(in == 657) begin
					state<=2;
					out<=51;
				end
				if(in == 658) begin
					state<=2;
					out<=52;
				end
				if(in == 659) begin
					state<=2;
					out<=53;
				end
				if(in == 660) begin
					state<=2;
					out<=54;
				end
				if(in == 661) begin
					state<=2;
					out<=55;
				end
				if(in == 662) begin
					state<=2;
					out<=56;
				end
				if(in == 663) begin
					state<=2;
					out<=57;
				end
				if(in == 664) begin
					state<=2;
					out<=58;
				end
				if(in == 665) begin
					state<=2;
					out<=59;
				end
				if(in == 666) begin
					state<=2;
					out<=60;
				end
				if(in == 667) begin
					state<=2;
					out<=61;
				end
				if(in == 668) begin
					state<=2;
					out<=62;
				end
				if(in == 669) begin
					state<=2;
					out<=63;
				end
				if(in == 670) begin
					state<=2;
					out<=64;
				end
				if(in == 671) begin
					state<=2;
					out<=65;
				end
				if(in == 672) begin
					state<=2;
					out<=66;
				end
				if(in == 673) begin
					state<=2;
					out<=67;
				end
				if(in == 674) begin
					state<=2;
					out<=68;
				end
				if(in == 675) begin
					state<=2;
					out<=69;
				end
				if(in == 676) begin
					state<=2;
					out<=70;
				end
				if(in == 677) begin
					state<=2;
					out<=71;
				end
				if(in == 678) begin
					state<=2;
					out<=72;
				end
				if(in == 679) begin
					state<=2;
					out<=73;
				end
				if(in == 680) begin
					state<=2;
					out<=74;
				end
				if(in == 681) begin
					state<=2;
					out<=75;
				end
				if(in == 682) begin
					state<=2;
					out<=76;
				end
				if(in == 683) begin
					state<=2;
					out<=77;
				end
				if(in == 684) begin
					state<=2;
					out<=78;
				end
				if(in == 685) begin
					state<=3;
					out<=79;
				end
				if(in == 686) begin
					state<=2;
					out<=80;
				end
				if(in == 687) begin
					state<=3;
					out<=81;
				end
				if(in == 688) begin
					state<=2;
					out<=82;
				end
				if(in == 689) begin
					state<=3;
					out<=83;
				end
				if(in == 690) begin
					state<=2;
					out<=84;
				end
				if(in == 691) begin
					state<=3;
					out<=85;
				end
				if(in == 692) begin
					state<=2;
					out<=86;
				end
				if(in == 693) begin
					state<=3;
					out<=87;
				end
				if(in == 694) begin
					state<=2;
					out<=88;
				end
				if(in == 695) begin
					state<=3;
					out<=89;
				end
				if(in == 696) begin
					state<=2;
					out<=90;
				end
				if(in == 697) begin
					state<=3;
					out<=91;
				end
				if(in == 698) begin
					state<=2;
					out<=92;
				end
				if(in == 699) begin
					state<=3;
					out<=93;
				end
				if(in == 700) begin
					state<=2;
					out<=94;
				end
				if(in == 701) begin
					state<=3;
					out<=95;
				end
				if(in == 702) begin
					state<=2;
					out<=96;
				end
				if(in == 703) begin
					state<=2;
					out<=97;
				end
				if(in == 704) begin
					state<=2;
					out<=98;
				end
				if(in == 705) begin
					state<=2;
					out<=99;
				end
				if(in == 706) begin
					state<=2;
					out<=100;
				end
				if(in == 707) begin
					state<=2;
					out<=101;
				end
				if(in == 708) begin
					state<=2;
					out<=102;
				end
				if(in == 709) begin
					state<=2;
					out<=103;
				end
				if(in == 710) begin
					state<=2;
					out<=104;
				end
				if(in == 711) begin
					state<=2;
					out<=105;
				end
				if(in == 712) begin
					state<=2;
					out<=106;
				end
				if(in == 713) begin
					state<=2;
					out<=107;
				end
				if(in == 714) begin
					state<=2;
					out<=108;
				end
				if(in == 715) begin
					state<=2;
					out<=109;
				end
				if(in == 716) begin
					state<=2;
					out<=110;
				end
				if(in == 717) begin
					state<=2;
					out<=111;
				end
				if(in == 718) begin
					state<=2;
					out<=112;
				end
				if(in == 719) begin
					state<=2;
					out<=113;
				end
				if(in == 720) begin
					state<=2;
					out<=114;
				end
				if(in == 721) begin
					state<=2;
					out<=115;
				end
				if(in == 722) begin
					state<=2;
					out<=116;
				end
				if(in == 723) begin
					state<=2;
					out<=117;
				end
				if(in == 724) begin
					state<=2;
					out<=118;
				end
				if(in == 725) begin
					state<=2;
					out<=119;
				end
				if(in == 726) begin
					state<=2;
					out<=120;
				end
				if(in == 727) begin
					state<=2;
					out<=121;
				end
				if(in == 728) begin
					state<=2;
					out<=122;
				end
				if(in == 729) begin
					state<=2;
					out<=123;
				end
				if(in == 730) begin
					state<=2;
					out<=124;
				end
				if(in == 731) begin
					state<=2;
					out<=125;
				end
				if(in == 732) begin
					state<=2;
					out<=126;
				end
				if(in == 733) begin
					state<=2;
					out<=127;
				end
				if(in == 734) begin
					state<=2;
					out<=128;
				end
				if(in == 735) begin
					state<=2;
					out<=129;
				end
				if(in == 736) begin
					state<=2;
					out<=130;
				end
				if(in == 737) begin
					state<=2;
					out<=131;
				end
				if(in == 738) begin
					state<=2;
					out<=132;
				end
				if(in == 739) begin
					state<=2;
					out<=133;
				end
				if(in == 740) begin
					state<=2;
					out<=134;
				end
				if(in == 741) begin
					state<=2;
					out<=135;
				end
				if(in == 742) begin
					state<=2;
					out<=136;
				end
				if(in == 743) begin
					state<=2;
					out<=137;
				end
				if(in == 744) begin
					state<=2;
					out<=138;
				end
				if(in == 745) begin
					state<=2;
					out<=139;
				end
				if(in == 746) begin
					state<=2;
					out<=140;
				end
				if(in == 747) begin
					state<=2;
					out<=141;
				end
				if(in == 748) begin
					state<=2;
					out<=142;
				end
				if(in == 749) begin
					state<=3;
					out<=143;
				end
				if(in == 750) begin
					state<=2;
					out<=144;
				end
				if(in == 751) begin
					state<=3;
					out<=145;
				end
				if(in == 752) begin
					state<=2;
					out<=146;
				end
				if(in == 753) begin
					state<=3;
					out<=147;
				end
				if(in == 754) begin
					state<=2;
					out<=148;
				end
				if(in == 755) begin
					state<=2;
					out<=149;
				end
				if(in == 756) begin
					state<=2;
					out<=150;
				end
				if(in == 757) begin
					state<=2;
					out<=151;
				end
				if(in == 758) begin
					state<=2;
					out<=152;
				end
				if(in == 759) begin
					state<=2;
					out<=153;
				end
				if(in == 760) begin
					state<=2;
					out<=154;
				end
				if(in == 761) begin
					state<=2;
					out<=155;
				end
				if(in == 762) begin
					state<=2;
					out<=156;
				end
				if(in == 763) begin
					state<=2;
					out<=157;
				end
				if(in == 764) begin
					state<=2;
					out<=158;
				end
				if(in == 765) begin
					state<=2;
					out<=159;
				end
				if(in == 766) begin
					state<=2;
					out<=160;
				end
				if(in == 767) begin
					state<=2;
					out<=161;
				end
				if(in == 768) begin
					state<=2;
					out<=162;
				end
				if(in == 769) begin
					state<=2;
					out<=163;
				end
				if(in == 770) begin
					state<=2;
					out<=164;
				end
				if(in == 771) begin
					state<=2;
					out<=165;
				end
				if(in == 772) begin
					state<=2;
					out<=166;
				end
				if(in == 773) begin
					state<=2;
					out<=167;
				end
				if(in == 774) begin
					state<=2;
					out<=168;
				end
				if(in == 775) begin
					state<=2;
					out<=169;
				end
				if(in == 776) begin
					state<=2;
					out<=170;
				end
				if(in == 777) begin
					state<=2;
					out<=171;
				end
				if(in == 778) begin
					state<=2;
					out<=172;
				end
				if(in == 779) begin
					state<=2;
					out<=173;
				end
				if(in == 780) begin
					state<=2;
					out<=174;
				end
				if(in == 781) begin
					state<=2;
					out<=175;
				end
				if(in == 782) begin
					state<=2;
					out<=176;
				end
				if(in == 783) begin
					state<=2;
					out<=177;
				end
				if(in == 784) begin
					state<=2;
					out<=178;
				end
				if(in == 785) begin
					state<=2;
					out<=179;
				end
				if(in == 786) begin
					state<=2;
					out<=180;
				end
				if(in == 787) begin
					state<=2;
					out<=181;
				end
				if(in == 788) begin
					state<=2;
					out<=182;
				end
				if(in == 789) begin
					state<=2;
					out<=183;
				end
				if(in == 790) begin
					state<=2;
					out<=184;
				end
				if(in == 791) begin
					state<=2;
					out<=185;
				end
				if(in == 792) begin
					state<=2;
					out<=186;
				end
				if(in == 793) begin
					state<=2;
					out<=187;
				end
				if(in == 794) begin
					state<=2;
					out<=188;
				end
				if(in == 795) begin
					state<=2;
					out<=189;
				end
				if(in == 796) begin
					state<=2;
					out<=190;
				end
				if(in == 797) begin
					state<=2;
					out<=191;
				end
				if(in == 798) begin
					state<=2;
					out<=192;
				end
				if(in == 799) begin
					state<=2;
					out<=193;
				end
				if(in == 800) begin
					state<=2;
					out<=194;
				end
				if(in == 801) begin
					state<=3;
					out<=195;
				end
				if(in == 802) begin
					state<=2;
					out<=196;
				end
				if(in == 803) begin
					state<=3;
					out<=197;
				end
				if(in == 804) begin
					state<=2;
					out<=198;
				end
				if(in == 805) begin
					state<=3;
					out<=199;
				end
				if(in == 806) begin
					state<=2;
					out<=200;
				end
				if(in == 807) begin
					state<=3;
					out<=201;
				end
				if(in == 808) begin
					state<=2;
					out<=202;
				end
				if(in == 809) begin
					state<=3;
					out<=203;
				end
				if(in == 810) begin
					state<=2;
					out<=204;
				end
				if(in == 811) begin
					state<=3;
					out<=205;
				end
				if(in == 812) begin
					state<=2;
					out<=206;
				end
				if(in == 813) begin
					state<=3;
					out<=207;
				end
				if(in == 814) begin
					state<=2;
					out<=208;
				end
				if(in == 815) begin
					state<=3;
					out<=209;
				end
				if(in == 816) begin
					state<=2;
					out<=210;
				end
				if(in == 817) begin
					state<=3;
					out<=211;
				end
				if(in == 818) begin
					state<=2;
					out<=212;
				end
				if(in == 819) begin
					state<=2;
					out<=213;
				end
				if(in == 820) begin
					state<=2;
					out<=214;
				end
				if(in == 821) begin
					state<=2;
					out<=215;
				end
				if(in == 822) begin
					state<=2;
					out<=216;
				end
				if(in == 823) begin
					state<=2;
					out<=217;
				end
				if(in == 824) begin
					state<=2;
					out<=218;
				end
				if(in == 825) begin
					state<=2;
					out<=219;
				end
				if(in == 826) begin
					state<=2;
					out<=220;
				end
				if(in == 827) begin
					state<=2;
					out<=221;
				end
				if(in == 828) begin
					state<=2;
					out<=222;
				end
				if(in == 829) begin
					state<=2;
					out<=223;
				end
				if(in == 830) begin
					state<=2;
					out<=224;
				end
				if(in == 831) begin
					state<=2;
					out<=225;
				end
				if(in == 832) begin
					state<=2;
					out<=226;
				end
				if(in == 833) begin
					state<=2;
					out<=227;
				end
				if(in == 834) begin
					state<=2;
					out<=228;
				end
				if(in == 835) begin
					state<=2;
					out<=229;
				end
				if(in == 836) begin
					state<=2;
					out<=230;
				end
				if(in == 837) begin
					state<=2;
					out<=231;
				end
				if(in == 838) begin
					state<=2;
					out<=232;
				end
				if(in == 839) begin
					state<=2;
					out<=233;
				end
				if(in == 840) begin
					state<=2;
					out<=234;
				end
				if(in == 841) begin
					state<=2;
					out<=235;
				end
				if(in == 842) begin
					state<=2;
					out<=236;
				end
				if(in == 843) begin
					state<=2;
					out<=237;
				end
				if(in == 844) begin
					state<=2;
					out<=238;
				end
				if(in == 845) begin
					state<=2;
					out<=239;
				end
				if(in == 846) begin
					state<=2;
					out<=240;
				end
				if(in == 847) begin
					state<=2;
					out<=241;
				end
				if(in == 848) begin
					state<=2;
					out<=242;
				end
				if(in == 849) begin
					state<=2;
					out<=243;
				end
				if(in == 850) begin
					state<=2;
					out<=244;
				end
				if(in == 851) begin
					state<=2;
					out<=245;
				end
				if(in == 852) begin
					state<=2;
					out<=246;
				end
				if(in == 853) begin
					state<=2;
					out<=247;
				end
				if(in == 854) begin
					state<=2;
					out<=248;
				end
				if(in == 855) begin
					state<=2;
					out<=249;
				end
				if(in == 856) begin
					state<=2;
					out<=250;
				end
				if(in == 857) begin
					state<=2;
					out<=251;
				end
				if(in == 858) begin
					state<=2;
					out<=252;
				end
				if(in == 859) begin
					state<=2;
					out<=253;
				end
				if(in == 860) begin
					state<=2;
					out<=254;
				end
				if(in == 861) begin
					state<=2;
					out<=255;
				end
				if(in == 862) begin
					state<=2;
					out<=0;
				end
				if(in == 863) begin
					state<=2;
					out<=1;
				end
				if(in == 864) begin
					state<=2;
					out<=2;
				end
				if(in == 865) begin
					state<=3;
					out<=3;
				end
				if(in == 866) begin
					state<=2;
					out<=4;
				end
				if(in == 867) begin
					state<=3;
					out<=5;
				end
				if(in == 868) begin
					state<=2;
					out<=6;
				end
				if(in == 869) begin
					state<=3;
					out<=7;
				end
				if(in == 870) begin
					state<=2;
					out<=8;
				end
				if(in == 871) begin
					state<=2;
					out<=9;
				end
				if(in == 872) begin
					state<=2;
					out<=10;
				end
				if(in == 873) begin
					state<=2;
					out<=11;
				end
				if(in == 874) begin
					state<=2;
					out<=12;
				end
				if(in == 875) begin
					state<=2;
					out<=13;
				end
				if(in == 876) begin
					state<=2;
					out<=14;
				end
				if(in == 877) begin
					state<=2;
					out<=15;
				end
				if(in == 878) begin
					state<=2;
					out<=16;
				end
				if(in == 879) begin
					state<=2;
					out<=17;
				end
				if(in == 880) begin
					state<=2;
					out<=18;
				end
				if(in == 881) begin
					state<=2;
					out<=19;
				end
				if(in == 882) begin
					state<=2;
					out<=20;
				end
				if(in == 883) begin
					state<=2;
					out<=21;
				end
				if(in == 884) begin
					state<=2;
					out<=22;
				end
				if(in == 885) begin
					state<=2;
					out<=23;
				end
				if(in == 886) begin
					state<=2;
					out<=24;
				end
				if(in == 887) begin
					state<=2;
					out<=25;
				end
				if(in == 888) begin
					state<=2;
					out<=26;
				end
				if(in == 889) begin
					state<=2;
					out<=27;
				end
				if(in == 890) begin
					state<=2;
					out<=28;
				end
				if(in == 891) begin
					state<=2;
					out<=29;
				end
				if(in == 892) begin
					state<=2;
					out<=30;
				end
				if(in == 893) begin
					state<=2;
					out<=31;
				end
				if(in == 894) begin
					state<=2;
					out<=32;
				end
				if(in == 895) begin
					state<=2;
					out<=33;
				end
				if(in == 896) begin
					state<=2;
					out<=34;
				end
				if(in == 897) begin
					state<=2;
					out<=35;
				end
				if(in == 898) begin
					state<=2;
					out<=36;
				end
				if(in == 899) begin
					state<=2;
					out<=37;
				end
				if(in == 900) begin
					state<=2;
					out<=38;
				end
				if(in == 901) begin
					state<=2;
					out<=39;
				end
				if(in == 902) begin
					state<=2;
					out<=40;
				end
				if(in == 903) begin
					state<=2;
					out<=41;
				end
				if(in == 904) begin
					state<=2;
					out<=42;
				end
				if(in == 905) begin
					state<=2;
					out<=43;
				end
				if(in == 906) begin
					state<=2;
					out<=44;
				end
				if(in == 907) begin
					state<=2;
					out<=45;
				end
				if(in == 908) begin
					state<=2;
					out<=46;
				end
				if(in == 909) begin
					state<=2;
					out<=47;
				end
				if(in == 910) begin
					state<=2;
					out<=48;
				end
				if(in == 911) begin
					state<=2;
					out<=49;
				end
				if(in == 912) begin
					state<=2;
					out<=50;
				end
				if(in == 913) begin
					state<=2;
					out<=51;
				end
				if(in == 914) begin
					state<=2;
					out<=52;
				end
				if(in == 915) begin
					state<=2;
					out<=53;
				end
				if(in == 916) begin
					state<=2;
					out<=54;
				end
				if(in == 917) begin
					state<=3;
					out<=55;
				end
				if(in == 918) begin
					state<=2;
					out<=56;
				end
				if(in == 919) begin
					state<=3;
					out<=57;
				end
				if(in == 920) begin
					state<=2;
					out<=58;
				end
				if(in == 921) begin
					state<=3;
					out<=59;
				end
				if(in == 922) begin
					state<=2;
					out<=60;
				end
				if(in == 923) begin
					state<=3;
					out<=61;
				end
				if(in == 924) begin
					state<=2;
					out<=62;
				end
				if(in == 925) begin
					state<=3;
					out<=63;
				end
				if(in == 926) begin
					state<=2;
					out<=64;
				end
				if(in == 927) begin
					state<=3;
					out<=65;
				end
				if(in == 928) begin
					state<=2;
					out<=66;
				end
			end
			3: begin
				if(in == 0) begin
					state<=3;
					out<=67;
				end
				if(in == 1) begin
					state<=1;
					out<=68;
				end
				if(in == 2) begin
					state<=3;
					out<=69;
				end
				if(in == 3) begin
					state<=5;
					out<=70;
				end
				if(in == 4) begin
					state<=5;
					out<=71;
				end
				if(in == 5) begin
					state<=4;
					out<=72;
				end
				if(in == 6) begin
					state<=4;
					out<=73;
				end
				if(in == 7) begin
					state<=5;
					out<=74;
				end
				if(in == 8) begin
					state<=4;
					out<=75;
				end
				if(in == 9) begin
					state<=5;
					out<=76;
				end
				if(in == 10) begin
					state<=4;
					out<=77;
				end
				if(in == 11) begin
					state<=5;
					out<=78;
				end
				if(in == 12) begin
					state<=4;
					out<=79;
				end
				if(in == 13) begin
					state<=5;
					out<=80;
				end
				if(in == 14) begin
					state<=4;
					out<=81;
				end
				if(in == 15) begin
					state<=5;
					out<=82;
				end
				if(in == 16) begin
					state<=4;
					out<=83;
				end
				if(in == 17) begin
					state<=5;
					out<=84;
				end
				if(in == 18) begin
					state<=4;
					out<=85;
				end
				if(in == 19) begin
					state<=5;
					out<=86;
				end
				if(in == 20) begin
					state<=4;
					out<=87;
				end
				if(in == 21) begin
					state<=5;
					out<=88;
				end
				if(in == 22) begin
					state<=4;
					out<=89;
				end
				if(in == 23) begin
					state<=5;
					out<=90;
				end
				if(in == 24) begin
					state<=4;
					out<=91;
				end
				if(in == 25) begin
					state<=5;
					out<=92;
				end
				if(in == 26) begin
					state<=4;
					out<=93;
				end
				if(in == 27) begin
					state<=5;
					out<=94;
				end
				if(in == 28) begin
					state<=4;
					out<=95;
				end
				if(in == 29) begin
					state<=5;
					out<=96;
				end
				if(in == 30) begin
					state<=4;
					out<=97;
				end
				if(in == 31) begin
					state<=5;
					out<=98;
				end
				if(in == 32) begin
					state<=4;
					out<=99;
				end
				if(in == 33) begin
					state<=5;
					out<=100;
				end
				if(in == 34) begin
					state<=4;
					out<=101;
				end
				if(in == 35) begin
					state<=5;
					out<=102;
				end
				if(in == 36) begin
					state<=4;
					out<=103;
				end
				if(in == 37) begin
					state<=5;
					out<=104;
				end
				if(in == 38) begin
					state<=4;
					out<=105;
				end
				if(in == 39) begin
					state<=5;
					out<=106;
				end
				if(in == 40) begin
					state<=4;
					out<=107;
				end
				if(in == 41) begin
					state<=5;
					out<=108;
				end
				if(in == 42) begin
					state<=4;
					out<=109;
				end
				if(in == 43) begin
					state<=5;
					out<=110;
				end
				if(in == 44) begin
					state<=4;
					out<=111;
				end
				if(in == 45) begin
					state<=5;
					out<=112;
				end
				if(in == 46) begin
					state<=4;
					out<=113;
				end
				if(in == 47) begin
					state<=5;
					out<=114;
				end
				if(in == 48) begin
					state<=4;
					out<=115;
				end
				if(in == 49) begin
					state<=5;
					out<=116;
				end
				if(in == 50) begin
					state<=4;
					out<=117;
				end
				if(in == 51) begin
					state<=5;
					out<=118;
				end
				if(in == 52) begin
					state<=4;
					out<=119;
				end
				if(in == 53) begin
					state<=3;
					out<=120;
				end
				if(in == 54) begin
					state<=3;
					out<=121;
				end
				if(in == 55) begin
					state<=5;
					out<=122;
				end
				if(in == 56) begin
					state<=5;
					out<=123;
				end
				if(in == 57) begin
					state<=4;
					out<=124;
				end
				if(in == 58) begin
					state<=4;
					out<=125;
				end
				if(in == 59) begin
					state<=5;
					out<=126;
				end
				if(in == 60) begin
					state<=4;
					out<=127;
				end
				if(in == 61) begin
					state<=5;
					out<=128;
				end
				if(in == 62) begin
					state<=4;
					out<=129;
				end
				if(in == 63) begin
					state<=5;
					out<=130;
				end
				if(in == 64) begin
					state<=4;
					out<=131;
				end
				if(in == 65) begin
					state<=5;
					out<=132;
				end
				if(in == 66) begin
					state<=4;
					out<=133;
				end
				if(in == 67) begin
					state<=5;
					out<=134;
				end
				if(in == 68) begin
					state<=4;
					out<=135;
				end
				if(in == 69) begin
					state<=5;
					out<=136;
				end
				if(in == 70) begin
					state<=4;
					out<=137;
				end
				if(in == 71) begin
					state<=5;
					out<=138;
				end
				if(in == 72) begin
					state<=4;
					out<=139;
				end
				if(in == 73) begin
					state<=5;
					out<=140;
				end
				if(in == 74) begin
					state<=4;
					out<=141;
				end
				if(in == 75) begin
					state<=5;
					out<=142;
				end
				if(in == 76) begin
					state<=4;
					out<=143;
				end
				if(in == 77) begin
					state<=5;
					out<=144;
				end
				if(in == 78) begin
					state<=4;
					out<=145;
				end
				if(in == 79) begin
					state<=5;
					out<=146;
				end
				if(in == 80) begin
					state<=4;
					out<=147;
				end
				if(in == 81) begin
					state<=5;
					out<=148;
				end
				if(in == 82) begin
					state<=4;
					out<=149;
				end
				if(in == 83) begin
					state<=5;
					out<=150;
				end
				if(in == 84) begin
					state<=4;
					out<=151;
				end
				if(in == 85) begin
					state<=5;
					out<=152;
				end
				if(in == 86) begin
					state<=4;
					out<=153;
				end
				if(in == 87) begin
					state<=5;
					out<=154;
				end
				if(in == 88) begin
					state<=4;
					out<=155;
				end
				if(in == 89) begin
					state<=5;
					out<=156;
				end
				if(in == 90) begin
					state<=4;
					out<=157;
				end
				if(in == 91) begin
					state<=5;
					out<=158;
				end
				if(in == 92) begin
					state<=4;
					out<=159;
				end
				if(in == 93) begin
					state<=5;
					out<=160;
				end
				if(in == 94) begin
					state<=4;
					out<=161;
				end
				if(in == 95) begin
					state<=5;
					out<=162;
				end
				if(in == 96) begin
					state<=4;
					out<=163;
				end
				if(in == 97) begin
					state<=5;
					out<=164;
				end
				if(in == 98) begin
					state<=4;
					out<=165;
				end
				if(in == 99) begin
					state<=5;
					out<=166;
				end
				if(in == 100) begin
					state<=4;
					out<=167;
				end
				if(in == 101) begin
					state<=5;
					out<=168;
				end
				if(in == 102) begin
					state<=4;
					out<=169;
				end
				if(in == 103) begin
					state<=5;
					out<=170;
				end
				if(in == 104) begin
					state<=4;
					out<=171;
				end
				if(in == 105) begin
					state<=3;
					out<=172;
				end
				if(in == 106) begin
					state<=3;
					out<=173;
				end
				if(in == 107) begin
					state<=5;
					out<=174;
				end
				if(in == 108) begin
					state<=5;
					out<=175;
				end
				if(in == 109) begin
					state<=4;
					out<=176;
				end
				if(in == 110) begin
					state<=4;
					out<=177;
				end
				if(in == 111) begin
					state<=3;
					out<=178;
				end
				if(in == 112) begin
					state<=3;
					out<=179;
				end
				if(in == 113) begin
					state<=5;
					out<=180;
				end
				if(in == 114) begin
					state<=5;
					out<=181;
				end
				if(in == 115) begin
					state<=4;
					out<=182;
				end
				if(in == 116) begin
					state<=4;
					out<=183;
				end
				if(in == 117) begin
					state<=3;
					out<=184;
				end
				if(in == 118) begin
					state<=3;
					out<=185;
				end
				if(in == 119) begin
					state<=5;
					out<=186;
				end
				if(in == 120) begin
					state<=5;
					out<=187;
				end
				if(in == 121) begin
					state<=4;
					out<=188;
				end
				if(in == 122) begin
					state<=4;
					out<=189;
				end
				if(in == 123) begin
					state<=5;
					out<=190;
				end
				if(in == 124) begin
					state<=4;
					out<=191;
				end
				if(in == 125) begin
					state<=5;
					out<=192;
				end
				if(in == 126) begin
					state<=4;
					out<=193;
				end
				if(in == 127) begin
					state<=5;
					out<=194;
				end
				if(in == 128) begin
					state<=4;
					out<=195;
				end
				if(in == 129) begin
					state<=5;
					out<=196;
				end
				if(in == 130) begin
					state<=4;
					out<=197;
				end
				if(in == 131) begin
					state<=5;
					out<=198;
				end
				if(in == 132) begin
					state<=4;
					out<=199;
				end
				if(in == 133) begin
					state<=5;
					out<=200;
				end
				if(in == 134) begin
					state<=4;
					out<=201;
				end
				if(in == 135) begin
					state<=5;
					out<=202;
				end
				if(in == 136) begin
					state<=4;
					out<=203;
				end
				if(in == 137) begin
					state<=5;
					out<=204;
				end
				if(in == 138) begin
					state<=4;
					out<=205;
				end
				if(in == 139) begin
					state<=5;
					out<=206;
				end
				if(in == 140) begin
					state<=4;
					out<=207;
				end
				if(in == 141) begin
					state<=5;
					out<=208;
				end
				if(in == 142) begin
					state<=4;
					out<=209;
				end
				if(in == 143) begin
					state<=5;
					out<=210;
				end
				if(in == 144) begin
					state<=4;
					out<=211;
				end
				if(in == 145) begin
					state<=5;
					out<=212;
				end
				if(in == 146) begin
					state<=4;
					out<=213;
				end
				if(in == 147) begin
					state<=5;
					out<=214;
				end
				if(in == 148) begin
					state<=4;
					out<=215;
				end
				if(in == 149) begin
					state<=5;
					out<=216;
				end
				if(in == 150) begin
					state<=4;
					out<=217;
				end
				if(in == 151) begin
					state<=5;
					out<=218;
				end
				if(in == 152) begin
					state<=4;
					out<=219;
				end
				if(in == 153) begin
					state<=5;
					out<=220;
				end
				if(in == 154) begin
					state<=4;
					out<=221;
				end
				if(in == 155) begin
					state<=5;
					out<=222;
				end
				if(in == 156) begin
					state<=4;
					out<=223;
				end
				if(in == 157) begin
					state<=5;
					out<=224;
				end
				if(in == 158) begin
					state<=4;
					out<=225;
				end
				if(in == 159) begin
					state<=5;
					out<=226;
				end
				if(in == 160) begin
					state<=4;
					out<=227;
				end
				if(in == 161) begin
					state<=5;
					out<=228;
				end
				if(in == 162) begin
					state<=4;
					out<=229;
				end
				if(in == 163) begin
					state<=5;
					out<=230;
				end
				if(in == 164) begin
					state<=4;
					out<=231;
				end
				if(in == 165) begin
					state<=5;
					out<=232;
				end
				if(in == 166) begin
					state<=4;
					out<=233;
				end
				if(in == 167) begin
					state<=5;
					out<=234;
				end
				if(in == 168) begin
					state<=4;
					out<=235;
				end
				if(in == 169) begin
					state<=3;
					out<=236;
				end
				if(in == 170) begin
					state<=3;
					out<=237;
				end
				if(in == 171) begin
					state<=5;
					out<=238;
				end
				if(in == 172) begin
					state<=5;
					out<=239;
				end
				if(in == 173) begin
					state<=4;
					out<=240;
				end
				if(in == 174) begin
					state<=4;
					out<=241;
				end
				if(in == 175) begin
					state<=5;
					out<=242;
				end
				if(in == 176) begin
					state<=4;
					out<=243;
				end
				if(in == 177) begin
					state<=5;
					out<=244;
				end
				if(in == 178) begin
					state<=4;
					out<=245;
				end
				if(in == 179) begin
					state<=5;
					out<=246;
				end
				if(in == 180) begin
					state<=4;
					out<=247;
				end
				if(in == 181) begin
					state<=5;
					out<=248;
				end
				if(in == 182) begin
					state<=4;
					out<=249;
				end
				if(in == 183) begin
					state<=5;
					out<=250;
				end
				if(in == 184) begin
					state<=4;
					out<=251;
				end
				if(in == 185) begin
					state<=5;
					out<=252;
				end
				if(in == 186) begin
					state<=4;
					out<=253;
				end
				if(in == 187) begin
					state<=5;
					out<=254;
				end
				if(in == 188) begin
					state<=4;
					out<=255;
				end
				if(in == 189) begin
					state<=5;
					out<=0;
				end
				if(in == 190) begin
					state<=4;
					out<=1;
				end
				if(in == 191) begin
					state<=5;
					out<=2;
				end
				if(in == 192) begin
					state<=4;
					out<=3;
				end
				if(in == 193) begin
					state<=5;
					out<=4;
				end
				if(in == 194) begin
					state<=4;
					out<=5;
				end
				if(in == 195) begin
					state<=5;
					out<=6;
				end
				if(in == 196) begin
					state<=4;
					out<=7;
				end
				if(in == 197) begin
					state<=5;
					out<=8;
				end
				if(in == 198) begin
					state<=4;
					out<=9;
				end
				if(in == 199) begin
					state<=5;
					out<=10;
				end
				if(in == 200) begin
					state<=4;
					out<=11;
				end
				if(in == 201) begin
					state<=5;
					out<=12;
				end
				if(in == 202) begin
					state<=4;
					out<=13;
				end
				if(in == 203) begin
					state<=5;
					out<=14;
				end
				if(in == 204) begin
					state<=4;
					out<=15;
				end
				if(in == 205) begin
					state<=5;
					out<=16;
				end
				if(in == 206) begin
					state<=4;
					out<=17;
				end
				if(in == 207) begin
					state<=5;
					out<=18;
				end
				if(in == 208) begin
					state<=4;
					out<=19;
				end
				if(in == 209) begin
					state<=5;
					out<=20;
				end
				if(in == 210) begin
					state<=4;
					out<=21;
				end
				if(in == 211) begin
					state<=5;
					out<=22;
				end
				if(in == 212) begin
					state<=4;
					out<=23;
				end
				if(in == 213) begin
					state<=5;
					out<=24;
				end
				if(in == 214) begin
					state<=4;
					out<=25;
				end
				if(in == 215) begin
					state<=5;
					out<=26;
				end
				if(in == 216) begin
					state<=4;
					out<=27;
				end
				if(in == 217) begin
					state<=5;
					out<=28;
				end
				if(in == 218) begin
					state<=4;
					out<=29;
				end
				if(in == 219) begin
					state<=5;
					out<=30;
				end
				if(in == 220) begin
					state<=4;
					out<=31;
				end
				if(in == 221) begin
					state<=3;
					out<=32;
				end
				if(in == 222) begin
					state<=3;
					out<=33;
				end
				if(in == 223) begin
					state<=5;
					out<=34;
				end
				if(in == 224) begin
					state<=5;
					out<=35;
				end
				if(in == 225) begin
					state<=4;
					out<=36;
				end
				if(in == 226) begin
					state<=4;
					out<=37;
				end
				if(in == 227) begin
					state<=3;
					out<=38;
				end
				if(in == 228) begin
					state<=3;
					out<=39;
				end
				if(in == 229) begin
					state<=5;
					out<=40;
				end
				if(in == 230) begin
					state<=5;
					out<=41;
				end
				if(in == 231) begin
					state<=4;
					out<=42;
				end
				if(in == 232) begin
					state<=4;
					out<=43;
				end
				if(in == 233) begin
					state<=3;
					out<=44;
				end
				if(in == 234) begin
					state<=3;
					out<=45;
				end
				if(in == 235) begin
					state<=5;
					out<=46;
				end
				if(in == 236) begin
					state<=5;
					out<=47;
				end
				if(in == 237) begin
					state<=4;
					out<=48;
				end
				if(in == 238) begin
					state<=4;
					out<=49;
				end
				if(in == 239) begin
					state<=5;
					out<=50;
				end
				if(in == 240) begin
					state<=4;
					out<=51;
				end
				if(in == 241) begin
					state<=5;
					out<=52;
				end
				if(in == 242) begin
					state<=4;
					out<=53;
				end
				if(in == 243) begin
					state<=5;
					out<=54;
				end
				if(in == 244) begin
					state<=4;
					out<=55;
				end
				if(in == 245) begin
					state<=5;
					out<=56;
				end
				if(in == 246) begin
					state<=4;
					out<=57;
				end
				if(in == 247) begin
					state<=5;
					out<=58;
				end
				if(in == 248) begin
					state<=4;
					out<=59;
				end
				if(in == 249) begin
					state<=5;
					out<=60;
				end
				if(in == 250) begin
					state<=4;
					out<=61;
				end
				if(in == 251) begin
					state<=5;
					out<=62;
				end
				if(in == 252) begin
					state<=4;
					out<=63;
				end
				if(in == 253) begin
					state<=5;
					out<=64;
				end
				if(in == 254) begin
					state<=4;
					out<=65;
				end
				if(in == 255) begin
					state<=5;
					out<=66;
				end
				if(in == 256) begin
					state<=4;
					out<=67;
				end
				if(in == 257) begin
					state<=5;
					out<=68;
				end
				if(in == 258) begin
					state<=4;
					out<=69;
				end
				if(in == 259) begin
					state<=5;
					out<=70;
				end
				if(in == 260) begin
					state<=4;
					out<=71;
				end
				if(in == 261) begin
					state<=5;
					out<=72;
				end
				if(in == 262) begin
					state<=4;
					out<=73;
				end
				if(in == 263) begin
					state<=5;
					out<=74;
				end
				if(in == 264) begin
					state<=4;
					out<=75;
				end
				if(in == 265) begin
					state<=5;
					out<=76;
				end
				if(in == 266) begin
					state<=4;
					out<=77;
				end
				if(in == 267) begin
					state<=5;
					out<=78;
				end
				if(in == 268) begin
					state<=4;
					out<=79;
				end
				if(in == 269) begin
					state<=5;
					out<=80;
				end
				if(in == 270) begin
					state<=4;
					out<=81;
				end
				if(in == 271) begin
					state<=5;
					out<=82;
				end
				if(in == 272) begin
					state<=4;
					out<=83;
				end
				if(in == 273) begin
					state<=5;
					out<=84;
				end
				if(in == 274) begin
					state<=4;
					out<=85;
				end
				if(in == 275) begin
					state<=5;
					out<=86;
				end
				if(in == 276) begin
					state<=4;
					out<=87;
				end
				if(in == 277) begin
					state<=5;
					out<=88;
				end
				if(in == 278) begin
					state<=4;
					out<=89;
				end
				if(in == 279) begin
					state<=5;
					out<=90;
				end
				if(in == 280) begin
					state<=4;
					out<=91;
				end
				if(in == 281) begin
					state<=5;
					out<=92;
				end
				if(in == 282) begin
					state<=4;
					out<=93;
				end
				if(in == 283) begin
					state<=5;
					out<=94;
				end
				if(in == 284) begin
					state<=4;
					out<=95;
				end
				if(in == 285) begin
					state<=3;
					out<=96;
				end
				if(in == 286) begin
					state<=3;
					out<=97;
				end
				if(in == 287) begin
					state<=5;
					out<=98;
				end
				if(in == 288) begin
					state<=5;
					out<=99;
				end
				if(in == 289) begin
					state<=4;
					out<=100;
				end
				if(in == 290) begin
					state<=4;
					out<=101;
				end
				if(in == 291) begin
					state<=5;
					out<=102;
				end
				if(in == 292) begin
					state<=4;
					out<=103;
				end
				if(in == 293) begin
					state<=5;
					out<=104;
				end
				if(in == 294) begin
					state<=4;
					out<=105;
				end
				if(in == 295) begin
					state<=5;
					out<=106;
				end
				if(in == 296) begin
					state<=4;
					out<=107;
				end
				if(in == 297) begin
					state<=5;
					out<=108;
				end
				if(in == 298) begin
					state<=4;
					out<=109;
				end
				if(in == 299) begin
					state<=5;
					out<=110;
				end
				if(in == 300) begin
					state<=4;
					out<=111;
				end
				if(in == 301) begin
					state<=5;
					out<=112;
				end
				if(in == 302) begin
					state<=4;
					out<=113;
				end
				if(in == 303) begin
					state<=5;
					out<=114;
				end
				if(in == 304) begin
					state<=4;
					out<=115;
				end
				if(in == 305) begin
					state<=5;
					out<=116;
				end
				if(in == 306) begin
					state<=4;
					out<=117;
				end
				if(in == 307) begin
					state<=5;
					out<=118;
				end
				if(in == 308) begin
					state<=4;
					out<=119;
				end
				if(in == 309) begin
					state<=5;
					out<=120;
				end
				if(in == 310) begin
					state<=4;
					out<=121;
				end
				if(in == 311) begin
					state<=5;
					out<=122;
				end
				if(in == 312) begin
					state<=4;
					out<=123;
				end
				if(in == 313) begin
					state<=5;
					out<=124;
				end
				if(in == 314) begin
					state<=4;
					out<=125;
				end
				if(in == 315) begin
					state<=5;
					out<=126;
				end
				if(in == 316) begin
					state<=4;
					out<=127;
				end
				if(in == 317) begin
					state<=5;
					out<=128;
				end
				if(in == 318) begin
					state<=4;
					out<=129;
				end
				if(in == 319) begin
					state<=5;
					out<=130;
				end
				if(in == 320) begin
					state<=4;
					out<=131;
				end
				if(in == 321) begin
					state<=5;
					out<=132;
				end
				if(in == 322) begin
					state<=4;
					out<=133;
				end
				if(in == 323) begin
					state<=5;
					out<=134;
				end
				if(in == 324) begin
					state<=4;
					out<=135;
				end
				if(in == 325) begin
					state<=5;
					out<=136;
				end
				if(in == 326) begin
					state<=4;
					out<=137;
				end
				if(in == 327) begin
					state<=5;
					out<=138;
				end
				if(in == 328) begin
					state<=4;
					out<=139;
				end
				if(in == 329) begin
					state<=5;
					out<=140;
				end
				if(in == 330) begin
					state<=4;
					out<=141;
				end
				if(in == 331) begin
					state<=5;
					out<=142;
				end
				if(in == 332) begin
					state<=4;
					out<=143;
				end
				if(in == 333) begin
					state<=5;
					out<=144;
				end
				if(in == 334) begin
					state<=4;
					out<=145;
				end
				if(in == 335) begin
					state<=5;
					out<=146;
				end
				if(in == 336) begin
					state<=4;
					out<=147;
				end
				if(in == 337) begin
					state<=3;
					out<=148;
				end
				if(in == 338) begin
					state<=3;
					out<=149;
				end
				if(in == 339) begin
					state<=5;
					out<=150;
				end
				if(in == 340) begin
					state<=5;
					out<=151;
				end
				if(in == 341) begin
					state<=4;
					out<=152;
				end
				if(in == 342) begin
					state<=4;
					out<=153;
				end
				if(in == 343) begin
					state<=3;
					out<=154;
				end
				if(in == 344) begin
					state<=3;
					out<=155;
				end
				if(in == 345) begin
					state<=5;
					out<=156;
				end
				if(in == 346) begin
					state<=5;
					out<=157;
				end
				if(in == 347) begin
					state<=4;
					out<=158;
				end
				if(in == 348) begin
					state<=4;
					out<=159;
				end
				if(in == 349) begin
					state<=3;
					out<=160;
				end
				if(in == 350) begin
					state<=3;
					out<=161;
				end
				if(in == 351) begin
					state<=5;
					out<=162;
				end
				if(in == 352) begin
					state<=5;
					out<=163;
				end
				if(in == 353) begin
					state<=4;
					out<=164;
				end
				if(in == 354) begin
					state<=4;
					out<=165;
				end
				if(in == 355) begin
					state<=5;
					out<=166;
				end
				if(in == 356) begin
					state<=4;
					out<=167;
				end
				if(in == 357) begin
					state<=5;
					out<=168;
				end
				if(in == 358) begin
					state<=4;
					out<=169;
				end
				if(in == 359) begin
					state<=5;
					out<=170;
				end
				if(in == 360) begin
					state<=4;
					out<=171;
				end
				if(in == 361) begin
					state<=5;
					out<=172;
				end
				if(in == 362) begin
					state<=4;
					out<=173;
				end
				if(in == 363) begin
					state<=5;
					out<=174;
				end
				if(in == 364) begin
					state<=4;
					out<=175;
				end
				if(in == 365) begin
					state<=5;
					out<=176;
				end
				if(in == 366) begin
					state<=4;
					out<=177;
				end
				if(in == 367) begin
					state<=5;
					out<=178;
				end
				if(in == 368) begin
					state<=4;
					out<=179;
				end
				if(in == 369) begin
					state<=5;
					out<=180;
				end
				if(in == 370) begin
					state<=4;
					out<=181;
				end
				if(in == 371) begin
					state<=5;
					out<=182;
				end
				if(in == 372) begin
					state<=4;
					out<=183;
				end
				if(in == 373) begin
					state<=5;
					out<=184;
				end
				if(in == 374) begin
					state<=4;
					out<=185;
				end
				if(in == 375) begin
					state<=5;
					out<=186;
				end
				if(in == 376) begin
					state<=4;
					out<=187;
				end
				if(in == 377) begin
					state<=5;
					out<=188;
				end
				if(in == 378) begin
					state<=4;
					out<=189;
				end
				if(in == 379) begin
					state<=5;
					out<=190;
				end
				if(in == 380) begin
					state<=4;
					out<=191;
				end
				if(in == 381) begin
					state<=5;
					out<=192;
				end
				if(in == 382) begin
					state<=4;
					out<=193;
				end
				if(in == 383) begin
					state<=5;
					out<=194;
				end
				if(in == 384) begin
					state<=4;
					out<=195;
				end
				if(in == 385) begin
					state<=5;
					out<=196;
				end
				if(in == 386) begin
					state<=4;
					out<=197;
				end
				if(in == 387) begin
					state<=5;
					out<=198;
				end
				if(in == 388) begin
					state<=4;
					out<=199;
				end
				if(in == 389) begin
					state<=5;
					out<=200;
				end
				if(in == 390) begin
					state<=4;
					out<=201;
				end
				if(in == 391) begin
					state<=5;
					out<=202;
				end
				if(in == 392) begin
					state<=4;
					out<=203;
				end
				if(in == 393) begin
					state<=5;
					out<=204;
				end
				if(in == 394) begin
					state<=4;
					out<=205;
				end
				if(in == 395) begin
					state<=5;
					out<=206;
				end
				if(in == 396) begin
					state<=4;
					out<=207;
				end
				if(in == 397) begin
					state<=5;
					out<=208;
				end
				if(in == 398) begin
					state<=4;
					out<=209;
				end
				if(in == 399) begin
					state<=5;
					out<=210;
				end
				if(in == 400) begin
					state<=4;
					out<=211;
				end
				if(in == 401) begin
					state<=3;
					out<=212;
				end
				if(in == 402) begin
					state<=3;
					out<=213;
				end
				if(in == 403) begin
					state<=5;
					out<=214;
				end
				if(in == 404) begin
					state<=5;
					out<=215;
				end
				if(in == 405) begin
					state<=4;
					out<=216;
				end
				if(in == 406) begin
					state<=4;
					out<=217;
				end
				if(in == 407) begin
					state<=5;
					out<=218;
				end
				if(in == 408) begin
					state<=4;
					out<=219;
				end
				if(in == 409) begin
					state<=5;
					out<=220;
				end
				if(in == 410) begin
					state<=4;
					out<=221;
				end
				if(in == 411) begin
					state<=5;
					out<=222;
				end
				if(in == 412) begin
					state<=4;
					out<=223;
				end
				if(in == 413) begin
					state<=5;
					out<=224;
				end
				if(in == 414) begin
					state<=4;
					out<=225;
				end
				if(in == 415) begin
					state<=5;
					out<=226;
				end
				if(in == 416) begin
					state<=4;
					out<=227;
				end
				if(in == 417) begin
					state<=5;
					out<=228;
				end
				if(in == 418) begin
					state<=4;
					out<=229;
				end
				if(in == 419) begin
					state<=5;
					out<=230;
				end
				if(in == 420) begin
					state<=4;
					out<=231;
				end
				if(in == 421) begin
					state<=5;
					out<=232;
				end
				if(in == 422) begin
					state<=4;
					out<=233;
				end
				if(in == 423) begin
					state<=5;
					out<=234;
				end
				if(in == 424) begin
					state<=4;
					out<=235;
				end
				if(in == 425) begin
					state<=5;
					out<=236;
				end
				if(in == 426) begin
					state<=4;
					out<=237;
				end
				if(in == 427) begin
					state<=5;
					out<=238;
				end
				if(in == 428) begin
					state<=4;
					out<=239;
				end
				if(in == 429) begin
					state<=5;
					out<=240;
				end
				if(in == 430) begin
					state<=4;
					out<=241;
				end
				if(in == 431) begin
					state<=5;
					out<=242;
				end
				if(in == 432) begin
					state<=4;
					out<=243;
				end
				if(in == 433) begin
					state<=5;
					out<=244;
				end
				if(in == 434) begin
					state<=4;
					out<=245;
				end
				if(in == 435) begin
					state<=5;
					out<=246;
				end
				if(in == 436) begin
					state<=4;
					out<=247;
				end
				if(in == 437) begin
					state<=5;
					out<=248;
				end
				if(in == 438) begin
					state<=4;
					out<=249;
				end
				if(in == 439) begin
					state<=5;
					out<=250;
				end
				if(in == 440) begin
					state<=4;
					out<=251;
				end
				if(in == 441) begin
					state<=5;
					out<=252;
				end
				if(in == 442) begin
					state<=4;
					out<=253;
				end
				if(in == 443) begin
					state<=5;
					out<=254;
				end
				if(in == 444) begin
					state<=4;
					out<=255;
				end
				if(in == 445) begin
					state<=5;
					out<=0;
				end
				if(in == 446) begin
					state<=4;
					out<=1;
				end
				if(in == 447) begin
					state<=5;
					out<=2;
				end
				if(in == 448) begin
					state<=4;
					out<=3;
				end
				if(in == 449) begin
					state<=5;
					out<=4;
				end
				if(in == 450) begin
					state<=4;
					out<=5;
				end
				if(in == 451) begin
					state<=5;
					out<=6;
				end
				if(in == 452) begin
					state<=4;
					out<=7;
				end
				if(in == 453) begin
					state<=3;
					out<=8;
				end
				if(in == 454) begin
					state<=3;
					out<=9;
				end
				if(in == 455) begin
					state<=5;
					out<=10;
				end
				if(in == 456) begin
					state<=5;
					out<=11;
				end
				if(in == 457) begin
					state<=4;
					out<=12;
				end
				if(in == 458) begin
					state<=4;
					out<=13;
				end
				if(in == 459) begin
					state<=3;
					out<=14;
				end
				if(in == 460) begin
					state<=3;
					out<=15;
				end
				if(in == 461) begin
					state<=5;
					out<=16;
				end
				if(in == 462) begin
					state<=5;
					out<=17;
				end
				if(in == 463) begin
					state<=4;
					out<=18;
				end
				if(in == 464) begin
					state<=4;
					out<=19;
				end
				if(in == 465) begin
					state<=3;
					out<=20;
				end
				if(in == 466) begin
					state<=3;
					out<=21;
				end
				if(in == 467) begin
					state<=5;
					out<=22;
				end
				if(in == 468) begin
					state<=5;
					out<=23;
				end
				if(in == 469) begin
					state<=4;
					out<=24;
				end
				if(in == 470) begin
					state<=4;
					out<=25;
				end
				if(in == 471) begin
					state<=5;
					out<=26;
				end
				if(in == 472) begin
					state<=4;
					out<=27;
				end
				if(in == 473) begin
					state<=5;
					out<=28;
				end
				if(in == 474) begin
					state<=4;
					out<=29;
				end
				if(in == 475) begin
					state<=5;
					out<=30;
				end
				if(in == 476) begin
					state<=4;
					out<=31;
				end
				if(in == 477) begin
					state<=5;
					out<=32;
				end
				if(in == 478) begin
					state<=4;
					out<=33;
				end
				if(in == 479) begin
					state<=5;
					out<=34;
				end
				if(in == 480) begin
					state<=4;
					out<=35;
				end
				if(in == 481) begin
					state<=5;
					out<=36;
				end
				if(in == 482) begin
					state<=4;
					out<=37;
				end
				if(in == 483) begin
					state<=5;
					out<=38;
				end
				if(in == 484) begin
					state<=4;
					out<=39;
				end
				if(in == 485) begin
					state<=5;
					out<=40;
				end
				if(in == 486) begin
					state<=4;
					out<=41;
				end
				if(in == 487) begin
					state<=5;
					out<=42;
				end
				if(in == 488) begin
					state<=4;
					out<=43;
				end
				if(in == 489) begin
					state<=5;
					out<=44;
				end
				if(in == 490) begin
					state<=4;
					out<=45;
				end
				if(in == 491) begin
					state<=5;
					out<=46;
				end
				if(in == 492) begin
					state<=4;
					out<=47;
				end
				if(in == 493) begin
					state<=5;
					out<=48;
				end
				if(in == 494) begin
					state<=4;
					out<=49;
				end
				if(in == 495) begin
					state<=5;
					out<=50;
				end
				if(in == 496) begin
					state<=4;
					out<=51;
				end
				if(in == 497) begin
					state<=5;
					out<=52;
				end
				if(in == 498) begin
					state<=4;
					out<=53;
				end
				if(in == 499) begin
					state<=5;
					out<=54;
				end
				if(in == 500) begin
					state<=4;
					out<=55;
				end
				if(in == 501) begin
					state<=5;
					out<=56;
				end
				if(in == 502) begin
					state<=4;
					out<=57;
				end
				if(in == 503) begin
					state<=5;
					out<=58;
				end
				if(in == 504) begin
					state<=4;
					out<=59;
				end
				if(in == 505) begin
					state<=5;
					out<=60;
				end
				if(in == 506) begin
					state<=4;
					out<=61;
				end
				if(in == 507) begin
					state<=5;
					out<=62;
				end
				if(in == 508) begin
					state<=4;
					out<=63;
				end
				if(in == 509) begin
					state<=5;
					out<=64;
				end
				if(in == 510) begin
					state<=4;
					out<=65;
				end
				if(in == 511) begin
					state<=5;
					out<=66;
				end
				if(in == 512) begin
					state<=4;
					out<=67;
				end
				if(in == 513) begin
					state<=5;
					out<=68;
				end
				if(in == 514) begin
					state<=4;
					out<=69;
				end
				if(in == 515) begin
					state<=5;
					out<=70;
				end
				if(in == 516) begin
					state<=4;
					out<=71;
				end
				if(in == 517) begin
					state<=3;
					out<=72;
				end
				if(in == 518) begin
					state<=3;
					out<=73;
				end
				if(in == 519) begin
					state<=5;
					out<=74;
				end
				if(in == 520) begin
					state<=5;
					out<=75;
				end
				if(in == 521) begin
					state<=4;
					out<=76;
				end
				if(in == 522) begin
					state<=4;
					out<=77;
				end
				if(in == 523) begin
					state<=5;
					out<=78;
				end
				if(in == 524) begin
					state<=4;
					out<=79;
				end
				if(in == 525) begin
					state<=5;
					out<=80;
				end
				if(in == 526) begin
					state<=4;
					out<=81;
				end
				if(in == 527) begin
					state<=5;
					out<=82;
				end
				if(in == 528) begin
					state<=4;
					out<=83;
				end
				if(in == 529) begin
					state<=5;
					out<=84;
				end
				if(in == 530) begin
					state<=4;
					out<=85;
				end
				if(in == 531) begin
					state<=5;
					out<=86;
				end
				if(in == 532) begin
					state<=4;
					out<=87;
				end
				if(in == 533) begin
					state<=5;
					out<=88;
				end
				if(in == 534) begin
					state<=4;
					out<=89;
				end
				if(in == 535) begin
					state<=5;
					out<=90;
				end
				if(in == 536) begin
					state<=4;
					out<=91;
				end
				if(in == 537) begin
					state<=5;
					out<=92;
				end
				if(in == 538) begin
					state<=4;
					out<=93;
				end
				if(in == 539) begin
					state<=5;
					out<=94;
				end
				if(in == 540) begin
					state<=4;
					out<=95;
				end
				if(in == 541) begin
					state<=5;
					out<=96;
				end
				if(in == 542) begin
					state<=4;
					out<=97;
				end
				if(in == 543) begin
					state<=5;
					out<=98;
				end
				if(in == 544) begin
					state<=4;
					out<=99;
				end
				if(in == 545) begin
					state<=5;
					out<=100;
				end
				if(in == 546) begin
					state<=4;
					out<=101;
				end
				if(in == 547) begin
					state<=5;
					out<=102;
				end
				if(in == 548) begin
					state<=4;
					out<=103;
				end
				if(in == 549) begin
					state<=5;
					out<=104;
				end
				if(in == 550) begin
					state<=4;
					out<=105;
				end
				if(in == 551) begin
					state<=5;
					out<=106;
				end
				if(in == 552) begin
					state<=4;
					out<=107;
				end
				if(in == 553) begin
					state<=5;
					out<=108;
				end
				if(in == 554) begin
					state<=4;
					out<=109;
				end
				if(in == 555) begin
					state<=5;
					out<=110;
				end
				if(in == 556) begin
					state<=4;
					out<=111;
				end
				if(in == 557) begin
					state<=5;
					out<=112;
				end
				if(in == 558) begin
					state<=4;
					out<=113;
				end
				if(in == 559) begin
					state<=5;
					out<=114;
				end
				if(in == 560) begin
					state<=4;
					out<=115;
				end
				if(in == 561) begin
					state<=5;
					out<=116;
				end
				if(in == 562) begin
					state<=4;
					out<=117;
				end
				if(in == 563) begin
					state<=5;
					out<=118;
				end
				if(in == 564) begin
					state<=4;
					out<=119;
				end
				if(in == 565) begin
					state<=5;
					out<=120;
				end
				if(in == 566) begin
					state<=4;
					out<=121;
				end
				if(in == 567) begin
					state<=5;
					out<=122;
				end
				if(in == 568) begin
					state<=4;
					out<=123;
				end
				if(in == 569) begin
					state<=3;
					out<=124;
				end
				if(in == 570) begin
					state<=3;
					out<=125;
				end
				if(in == 571) begin
					state<=5;
					out<=126;
				end
				if(in == 572) begin
					state<=5;
					out<=127;
				end
				if(in == 573) begin
					state<=4;
					out<=128;
				end
				if(in == 574) begin
					state<=4;
					out<=129;
				end
				if(in == 575) begin
					state<=3;
					out<=130;
				end
				if(in == 576) begin
					state<=3;
					out<=131;
				end
				if(in == 577) begin
					state<=5;
					out<=132;
				end
				if(in == 578) begin
					state<=5;
					out<=133;
				end
				if(in == 579) begin
					state<=4;
					out<=134;
				end
				if(in == 580) begin
					state<=4;
					out<=135;
				end
				if(in == 581) begin
					state<=3;
					out<=136;
				end
				if(in == 582) begin
					state<=3;
					out<=137;
				end
				if(in == 583) begin
					state<=5;
					out<=138;
				end
				if(in == 584) begin
					state<=5;
					out<=139;
				end
				if(in == 585) begin
					state<=4;
					out<=140;
				end
				if(in == 586) begin
					state<=4;
					out<=141;
				end
				if(in == 587) begin
					state<=5;
					out<=142;
				end
				if(in == 588) begin
					state<=4;
					out<=143;
				end
				if(in == 589) begin
					state<=5;
					out<=144;
				end
				if(in == 590) begin
					state<=4;
					out<=145;
				end
				if(in == 591) begin
					state<=5;
					out<=146;
				end
				if(in == 592) begin
					state<=4;
					out<=147;
				end
				if(in == 593) begin
					state<=5;
					out<=148;
				end
				if(in == 594) begin
					state<=4;
					out<=149;
				end
				if(in == 595) begin
					state<=5;
					out<=150;
				end
				if(in == 596) begin
					state<=4;
					out<=151;
				end
				if(in == 597) begin
					state<=5;
					out<=152;
				end
				if(in == 598) begin
					state<=4;
					out<=153;
				end
				if(in == 599) begin
					state<=5;
					out<=154;
				end
				if(in == 600) begin
					state<=4;
					out<=155;
				end
				if(in == 601) begin
					state<=5;
					out<=156;
				end
				if(in == 602) begin
					state<=4;
					out<=157;
				end
				if(in == 603) begin
					state<=5;
					out<=158;
				end
				if(in == 604) begin
					state<=4;
					out<=159;
				end
				if(in == 605) begin
					state<=5;
					out<=160;
				end
				if(in == 606) begin
					state<=4;
					out<=161;
				end
				if(in == 607) begin
					state<=5;
					out<=162;
				end
				if(in == 608) begin
					state<=4;
					out<=163;
				end
				if(in == 609) begin
					state<=5;
					out<=164;
				end
				if(in == 610) begin
					state<=4;
					out<=165;
				end
				if(in == 611) begin
					state<=5;
					out<=166;
				end
				if(in == 612) begin
					state<=4;
					out<=167;
				end
				if(in == 613) begin
					state<=5;
					out<=168;
				end
				if(in == 614) begin
					state<=4;
					out<=169;
				end
				if(in == 615) begin
					state<=5;
					out<=170;
				end
				if(in == 616) begin
					state<=4;
					out<=171;
				end
				if(in == 617) begin
					state<=5;
					out<=172;
				end
				if(in == 618) begin
					state<=4;
					out<=173;
				end
				if(in == 619) begin
					state<=5;
					out<=174;
				end
				if(in == 620) begin
					state<=4;
					out<=175;
				end
				if(in == 621) begin
					state<=5;
					out<=176;
				end
				if(in == 622) begin
					state<=4;
					out<=177;
				end
				if(in == 623) begin
					state<=5;
					out<=178;
				end
				if(in == 624) begin
					state<=4;
					out<=179;
				end
				if(in == 625) begin
					state<=5;
					out<=180;
				end
				if(in == 626) begin
					state<=4;
					out<=181;
				end
				if(in == 627) begin
					state<=5;
					out<=182;
				end
				if(in == 628) begin
					state<=4;
					out<=183;
				end
				if(in == 629) begin
					state<=5;
					out<=184;
				end
				if(in == 630) begin
					state<=4;
					out<=185;
				end
				if(in == 631) begin
					state<=5;
					out<=186;
				end
				if(in == 632) begin
					state<=4;
					out<=187;
				end
				if(in == 633) begin
					state<=3;
					out<=188;
				end
				if(in == 634) begin
					state<=3;
					out<=189;
				end
				if(in == 635) begin
					state<=5;
					out<=190;
				end
				if(in == 636) begin
					state<=5;
					out<=191;
				end
				if(in == 637) begin
					state<=4;
					out<=192;
				end
				if(in == 638) begin
					state<=4;
					out<=193;
				end
				if(in == 639) begin
					state<=5;
					out<=194;
				end
				if(in == 640) begin
					state<=4;
					out<=195;
				end
				if(in == 641) begin
					state<=5;
					out<=196;
				end
				if(in == 642) begin
					state<=4;
					out<=197;
				end
				if(in == 643) begin
					state<=5;
					out<=198;
				end
				if(in == 644) begin
					state<=4;
					out<=199;
				end
				if(in == 645) begin
					state<=5;
					out<=200;
				end
				if(in == 646) begin
					state<=4;
					out<=201;
				end
				if(in == 647) begin
					state<=5;
					out<=202;
				end
				if(in == 648) begin
					state<=4;
					out<=203;
				end
				if(in == 649) begin
					state<=5;
					out<=204;
				end
				if(in == 650) begin
					state<=4;
					out<=205;
				end
				if(in == 651) begin
					state<=5;
					out<=206;
				end
				if(in == 652) begin
					state<=4;
					out<=207;
				end
				if(in == 653) begin
					state<=5;
					out<=208;
				end
				if(in == 654) begin
					state<=4;
					out<=209;
				end
				if(in == 655) begin
					state<=5;
					out<=210;
				end
				if(in == 656) begin
					state<=4;
					out<=211;
				end
				if(in == 657) begin
					state<=5;
					out<=212;
				end
				if(in == 658) begin
					state<=4;
					out<=213;
				end
				if(in == 659) begin
					state<=5;
					out<=214;
				end
				if(in == 660) begin
					state<=4;
					out<=215;
				end
				if(in == 661) begin
					state<=5;
					out<=216;
				end
				if(in == 662) begin
					state<=4;
					out<=217;
				end
				if(in == 663) begin
					state<=5;
					out<=218;
				end
				if(in == 664) begin
					state<=4;
					out<=219;
				end
				if(in == 665) begin
					state<=5;
					out<=220;
				end
				if(in == 666) begin
					state<=4;
					out<=221;
				end
				if(in == 667) begin
					state<=5;
					out<=222;
				end
				if(in == 668) begin
					state<=4;
					out<=223;
				end
				if(in == 669) begin
					state<=5;
					out<=224;
				end
				if(in == 670) begin
					state<=4;
					out<=225;
				end
				if(in == 671) begin
					state<=5;
					out<=226;
				end
				if(in == 672) begin
					state<=4;
					out<=227;
				end
				if(in == 673) begin
					state<=5;
					out<=228;
				end
				if(in == 674) begin
					state<=4;
					out<=229;
				end
				if(in == 675) begin
					state<=5;
					out<=230;
				end
				if(in == 676) begin
					state<=4;
					out<=231;
				end
				if(in == 677) begin
					state<=5;
					out<=232;
				end
				if(in == 678) begin
					state<=4;
					out<=233;
				end
				if(in == 679) begin
					state<=5;
					out<=234;
				end
				if(in == 680) begin
					state<=4;
					out<=235;
				end
				if(in == 681) begin
					state<=5;
					out<=236;
				end
				if(in == 682) begin
					state<=4;
					out<=237;
				end
				if(in == 683) begin
					state<=5;
					out<=238;
				end
				if(in == 684) begin
					state<=4;
					out<=239;
				end
				if(in == 685) begin
					state<=3;
					out<=240;
				end
				if(in == 686) begin
					state<=3;
					out<=241;
				end
				if(in == 687) begin
					state<=5;
					out<=242;
				end
				if(in == 688) begin
					state<=5;
					out<=243;
				end
				if(in == 689) begin
					state<=4;
					out<=244;
				end
				if(in == 690) begin
					state<=4;
					out<=245;
				end
				if(in == 691) begin
					state<=3;
					out<=246;
				end
				if(in == 692) begin
					state<=3;
					out<=247;
				end
				if(in == 693) begin
					state<=5;
					out<=248;
				end
				if(in == 694) begin
					state<=5;
					out<=249;
				end
				if(in == 695) begin
					state<=4;
					out<=250;
				end
				if(in == 696) begin
					state<=4;
					out<=251;
				end
				if(in == 697) begin
					state<=3;
					out<=252;
				end
				if(in == 698) begin
					state<=3;
					out<=253;
				end
				if(in == 699) begin
					state<=5;
					out<=254;
				end
				if(in == 700) begin
					state<=5;
					out<=255;
				end
				if(in == 701) begin
					state<=4;
					out<=0;
				end
				if(in == 702) begin
					state<=4;
					out<=1;
				end
				if(in == 703) begin
					state<=5;
					out<=2;
				end
				if(in == 704) begin
					state<=4;
					out<=3;
				end
				if(in == 705) begin
					state<=5;
					out<=4;
				end
				if(in == 706) begin
					state<=4;
					out<=5;
				end
				if(in == 707) begin
					state<=5;
					out<=6;
				end
				if(in == 708) begin
					state<=4;
					out<=7;
				end
				if(in == 709) begin
					state<=5;
					out<=8;
				end
				if(in == 710) begin
					state<=4;
					out<=9;
				end
				if(in == 711) begin
					state<=5;
					out<=10;
				end
				if(in == 712) begin
					state<=4;
					out<=11;
				end
				if(in == 713) begin
					state<=5;
					out<=12;
				end
				if(in == 714) begin
					state<=4;
					out<=13;
				end
				if(in == 715) begin
					state<=5;
					out<=14;
				end
				if(in == 716) begin
					state<=4;
					out<=15;
				end
				if(in == 717) begin
					state<=5;
					out<=16;
				end
				if(in == 718) begin
					state<=4;
					out<=17;
				end
				if(in == 719) begin
					state<=5;
					out<=18;
				end
				if(in == 720) begin
					state<=4;
					out<=19;
				end
				if(in == 721) begin
					state<=5;
					out<=20;
				end
				if(in == 722) begin
					state<=4;
					out<=21;
				end
				if(in == 723) begin
					state<=5;
					out<=22;
				end
				if(in == 724) begin
					state<=4;
					out<=23;
				end
				if(in == 725) begin
					state<=5;
					out<=24;
				end
				if(in == 726) begin
					state<=4;
					out<=25;
				end
				if(in == 727) begin
					state<=5;
					out<=26;
				end
				if(in == 728) begin
					state<=4;
					out<=27;
				end
				if(in == 729) begin
					state<=5;
					out<=28;
				end
				if(in == 730) begin
					state<=4;
					out<=29;
				end
				if(in == 731) begin
					state<=5;
					out<=30;
				end
				if(in == 732) begin
					state<=4;
					out<=31;
				end
				if(in == 733) begin
					state<=5;
					out<=32;
				end
				if(in == 734) begin
					state<=4;
					out<=33;
				end
				if(in == 735) begin
					state<=5;
					out<=34;
				end
				if(in == 736) begin
					state<=4;
					out<=35;
				end
				if(in == 737) begin
					state<=5;
					out<=36;
				end
				if(in == 738) begin
					state<=4;
					out<=37;
				end
				if(in == 739) begin
					state<=5;
					out<=38;
				end
				if(in == 740) begin
					state<=4;
					out<=39;
				end
				if(in == 741) begin
					state<=5;
					out<=40;
				end
				if(in == 742) begin
					state<=4;
					out<=41;
				end
				if(in == 743) begin
					state<=5;
					out<=42;
				end
				if(in == 744) begin
					state<=4;
					out<=43;
				end
				if(in == 745) begin
					state<=5;
					out<=44;
				end
				if(in == 746) begin
					state<=4;
					out<=45;
				end
				if(in == 747) begin
					state<=5;
					out<=46;
				end
				if(in == 748) begin
					state<=4;
					out<=47;
				end
				if(in == 749) begin
					state<=3;
					out<=48;
				end
				if(in == 750) begin
					state<=3;
					out<=49;
				end
				if(in == 751) begin
					state<=5;
					out<=50;
				end
				if(in == 752) begin
					state<=5;
					out<=51;
				end
				if(in == 753) begin
					state<=4;
					out<=52;
				end
				if(in == 754) begin
					state<=4;
					out<=53;
				end
				if(in == 755) begin
					state<=5;
					out<=54;
				end
				if(in == 756) begin
					state<=4;
					out<=55;
				end
				if(in == 757) begin
					state<=5;
					out<=56;
				end
				if(in == 758) begin
					state<=4;
					out<=57;
				end
				if(in == 759) begin
					state<=5;
					out<=58;
				end
				if(in == 760) begin
					state<=4;
					out<=59;
				end
				if(in == 761) begin
					state<=5;
					out<=60;
				end
				if(in == 762) begin
					state<=4;
					out<=61;
				end
				if(in == 763) begin
					state<=5;
					out<=62;
				end
				if(in == 764) begin
					state<=4;
					out<=63;
				end
				if(in == 765) begin
					state<=5;
					out<=64;
				end
				if(in == 766) begin
					state<=4;
					out<=65;
				end
				if(in == 767) begin
					state<=5;
					out<=66;
				end
				if(in == 768) begin
					state<=4;
					out<=67;
				end
				if(in == 769) begin
					state<=5;
					out<=68;
				end
				if(in == 770) begin
					state<=4;
					out<=69;
				end
				if(in == 771) begin
					state<=5;
					out<=70;
				end
				if(in == 772) begin
					state<=4;
					out<=71;
				end
				if(in == 773) begin
					state<=5;
					out<=72;
				end
				if(in == 774) begin
					state<=4;
					out<=73;
				end
				if(in == 775) begin
					state<=5;
					out<=74;
				end
				if(in == 776) begin
					state<=4;
					out<=75;
				end
				if(in == 777) begin
					state<=5;
					out<=76;
				end
				if(in == 778) begin
					state<=4;
					out<=77;
				end
				if(in == 779) begin
					state<=5;
					out<=78;
				end
				if(in == 780) begin
					state<=4;
					out<=79;
				end
				if(in == 781) begin
					state<=5;
					out<=80;
				end
				if(in == 782) begin
					state<=4;
					out<=81;
				end
				if(in == 783) begin
					state<=5;
					out<=82;
				end
				if(in == 784) begin
					state<=4;
					out<=83;
				end
				if(in == 785) begin
					state<=5;
					out<=84;
				end
				if(in == 786) begin
					state<=4;
					out<=85;
				end
				if(in == 787) begin
					state<=5;
					out<=86;
				end
				if(in == 788) begin
					state<=4;
					out<=87;
				end
				if(in == 789) begin
					state<=5;
					out<=88;
				end
				if(in == 790) begin
					state<=4;
					out<=89;
				end
				if(in == 791) begin
					state<=5;
					out<=90;
				end
				if(in == 792) begin
					state<=4;
					out<=91;
				end
				if(in == 793) begin
					state<=5;
					out<=92;
				end
				if(in == 794) begin
					state<=4;
					out<=93;
				end
				if(in == 795) begin
					state<=5;
					out<=94;
				end
				if(in == 796) begin
					state<=4;
					out<=95;
				end
				if(in == 797) begin
					state<=5;
					out<=96;
				end
				if(in == 798) begin
					state<=4;
					out<=97;
				end
				if(in == 799) begin
					state<=5;
					out<=98;
				end
				if(in == 800) begin
					state<=4;
					out<=99;
				end
				if(in == 801) begin
					state<=3;
					out<=100;
				end
				if(in == 802) begin
					state<=3;
					out<=101;
				end
				if(in == 803) begin
					state<=5;
					out<=102;
				end
				if(in == 804) begin
					state<=5;
					out<=103;
				end
				if(in == 805) begin
					state<=4;
					out<=104;
				end
				if(in == 806) begin
					state<=4;
					out<=105;
				end
				if(in == 807) begin
					state<=3;
					out<=106;
				end
				if(in == 808) begin
					state<=3;
					out<=107;
				end
				if(in == 809) begin
					state<=5;
					out<=108;
				end
				if(in == 810) begin
					state<=5;
					out<=109;
				end
				if(in == 811) begin
					state<=4;
					out<=110;
				end
				if(in == 812) begin
					state<=4;
					out<=111;
				end
				if(in == 813) begin
					state<=3;
					out<=112;
				end
				if(in == 814) begin
					state<=3;
					out<=113;
				end
				if(in == 815) begin
					state<=5;
					out<=114;
				end
				if(in == 816) begin
					state<=5;
					out<=115;
				end
				if(in == 817) begin
					state<=4;
					out<=116;
				end
				if(in == 818) begin
					state<=4;
					out<=117;
				end
				if(in == 819) begin
					state<=5;
					out<=118;
				end
				if(in == 820) begin
					state<=4;
					out<=119;
				end
				if(in == 821) begin
					state<=5;
					out<=120;
				end
				if(in == 822) begin
					state<=4;
					out<=121;
				end
				if(in == 823) begin
					state<=5;
					out<=122;
				end
				if(in == 824) begin
					state<=4;
					out<=123;
				end
				if(in == 825) begin
					state<=5;
					out<=124;
				end
				if(in == 826) begin
					state<=4;
					out<=125;
				end
				if(in == 827) begin
					state<=5;
					out<=126;
				end
				if(in == 828) begin
					state<=4;
					out<=127;
				end
				if(in == 829) begin
					state<=5;
					out<=128;
				end
				if(in == 830) begin
					state<=4;
					out<=129;
				end
				if(in == 831) begin
					state<=5;
					out<=130;
				end
				if(in == 832) begin
					state<=4;
					out<=131;
				end
				if(in == 833) begin
					state<=5;
					out<=132;
				end
				if(in == 834) begin
					state<=4;
					out<=133;
				end
				if(in == 835) begin
					state<=5;
					out<=134;
				end
				if(in == 836) begin
					state<=4;
					out<=135;
				end
				if(in == 837) begin
					state<=5;
					out<=136;
				end
				if(in == 838) begin
					state<=4;
					out<=137;
				end
				if(in == 839) begin
					state<=5;
					out<=138;
				end
				if(in == 840) begin
					state<=4;
					out<=139;
				end
				if(in == 841) begin
					state<=5;
					out<=140;
				end
				if(in == 842) begin
					state<=4;
					out<=141;
				end
				if(in == 843) begin
					state<=5;
					out<=142;
				end
				if(in == 844) begin
					state<=4;
					out<=143;
				end
				if(in == 845) begin
					state<=5;
					out<=144;
				end
				if(in == 846) begin
					state<=4;
					out<=145;
				end
				if(in == 847) begin
					state<=5;
					out<=146;
				end
				if(in == 848) begin
					state<=4;
					out<=147;
				end
				if(in == 849) begin
					state<=5;
					out<=148;
				end
				if(in == 850) begin
					state<=4;
					out<=149;
				end
				if(in == 851) begin
					state<=5;
					out<=150;
				end
				if(in == 852) begin
					state<=4;
					out<=151;
				end
				if(in == 853) begin
					state<=5;
					out<=152;
				end
				if(in == 854) begin
					state<=4;
					out<=153;
				end
				if(in == 855) begin
					state<=5;
					out<=154;
				end
				if(in == 856) begin
					state<=4;
					out<=155;
				end
				if(in == 857) begin
					state<=5;
					out<=156;
				end
				if(in == 858) begin
					state<=4;
					out<=157;
				end
				if(in == 859) begin
					state<=5;
					out<=158;
				end
				if(in == 860) begin
					state<=4;
					out<=159;
				end
				if(in == 861) begin
					state<=5;
					out<=160;
				end
				if(in == 862) begin
					state<=4;
					out<=161;
				end
				if(in == 863) begin
					state<=5;
					out<=162;
				end
				if(in == 864) begin
					state<=4;
					out<=163;
				end
				if(in == 865) begin
					state<=3;
					out<=164;
				end
				if(in == 866) begin
					state<=3;
					out<=165;
				end
				if(in == 867) begin
					state<=5;
					out<=166;
				end
				if(in == 868) begin
					state<=5;
					out<=167;
				end
				if(in == 869) begin
					state<=4;
					out<=168;
				end
				if(in == 870) begin
					state<=4;
					out<=169;
				end
				if(in == 871) begin
					state<=5;
					out<=170;
				end
				if(in == 872) begin
					state<=4;
					out<=171;
				end
				if(in == 873) begin
					state<=5;
					out<=172;
				end
				if(in == 874) begin
					state<=4;
					out<=173;
				end
				if(in == 875) begin
					state<=5;
					out<=174;
				end
				if(in == 876) begin
					state<=4;
					out<=175;
				end
				if(in == 877) begin
					state<=5;
					out<=176;
				end
				if(in == 878) begin
					state<=4;
					out<=177;
				end
				if(in == 879) begin
					state<=5;
					out<=178;
				end
				if(in == 880) begin
					state<=4;
					out<=179;
				end
				if(in == 881) begin
					state<=5;
					out<=180;
				end
				if(in == 882) begin
					state<=4;
					out<=181;
				end
				if(in == 883) begin
					state<=5;
					out<=182;
				end
				if(in == 884) begin
					state<=4;
					out<=183;
				end
				if(in == 885) begin
					state<=5;
					out<=184;
				end
				if(in == 886) begin
					state<=4;
					out<=185;
				end
				if(in == 887) begin
					state<=5;
					out<=186;
				end
				if(in == 888) begin
					state<=4;
					out<=187;
				end
				if(in == 889) begin
					state<=5;
					out<=188;
				end
				if(in == 890) begin
					state<=4;
					out<=189;
				end
				if(in == 891) begin
					state<=5;
					out<=190;
				end
				if(in == 892) begin
					state<=4;
					out<=191;
				end
				if(in == 893) begin
					state<=5;
					out<=192;
				end
				if(in == 894) begin
					state<=4;
					out<=193;
				end
				if(in == 895) begin
					state<=5;
					out<=194;
				end
				if(in == 896) begin
					state<=4;
					out<=195;
				end
				if(in == 897) begin
					state<=5;
					out<=196;
				end
				if(in == 898) begin
					state<=4;
					out<=197;
				end
				if(in == 899) begin
					state<=5;
					out<=198;
				end
				if(in == 900) begin
					state<=4;
					out<=199;
				end
				if(in == 901) begin
					state<=5;
					out<=200;
				end
				if(in == 902) begin
					state<=4;
					out<=201;
				end
				if(in == 903) begin
					state<=5;
					out<=202;
				end
				if(in == 904) begin
					state<=4;
					out<=203;
				end
				if(in == 905) begin
					state<=5;
					out<=204;
				end
				if(in == 906) begin
					state<=4;
					out<=205;
				end
				if(in == 907) begin
					state<=5;
					out<=206;
				end
				if(in == 908) begin
					state<=4;
					out<=207;
				end
				if(in == 909) begin
					state<=5;
					out<=208;
				end
				if(in == 910) begin
					state<=4;
					out<=209;
				end
				if(in == 911) begin
					state<=5;
					out<=210;
				end
				if(in == 912) begin
					state<=4;
					out<=211;
				end
				if(in == 913) begin
					state<=5;
					out<=212;
				end
				if(in == 914) begin
					state<=4;
					out<=213;
				end
				if(in == 915) begin
					state<=5;
					out<=214;
				end
				if(in == 916) begin
					state<=4;
					out<=215;
				end
				if(in == 917) begin
					state<=3;
					out<=216;
				end
				if(in == 918) begin
					state<=3;
					out<=217;
				end
				if(in == 919) begin
					state<=5;
					out<=218;
				end
				if(in == 920) begin
					state<=5;
					out<=219;
				end
				if(in == 921) begin
					state<=4;
					out<=220;
				end
				if(in == 922) begin
					state<=4;
					out<=221;
				end
				if(in == 923) begin
					state<=3;
					out<=222;
				end
				if(in == 924) begin
					state<=3;
					out<=223;
				end
				if(in == 925) begin
					state<=5;
					out<=224;
				end
				if(in == 926) begin
					state<=5;
					out<=225;
				end
				if(in == 927) begin
					state<=4;
					out<=226;
				end
				if(in == 928) begin
					state<=4;
					out<=227;
				end
			end
			4: begin
				if(in == 0) begin
					state<=3;
					out<=228;
				end
				if(in == 1) begin
					state<=1;
					out<=229;
				end
				if(in == 2) begin
					state<=4;
					out<=230;
				end
				if(in == 3) begin
					state<=3;
					out<=231;
				end
				if(in == 4) begin
					state<=5;
					out<=232;
				end
				if(in == 5) begin
					state<=3;
					out<=233;
				end
				if(in == 6) begin
					state<=5;
					out<=234;
				end
				if(in == 7) begin
					state<=5;
					out<=235;
				end
				if(in == 8) begin
					state<=5;
					out<=236;
				end
				if(in == 9) begin
					state<=5;
					out<=237;
				end
				if(in == 10) begin
					state<=5;
					out<=238;
				end
				if(in == 11) begin
					state<=5;
					out<=239;
				end
				if(in == 12) begin
					state<=5;
					out<=240;
				end
				if(in == 13) begin
					state<=5;
					out<=241;
				end
				if(in == 14) begin
					state<=5;
					out<=242;
				end
				if(in == 15) begin
					state<=5;
					out<=243;
				end
				if(in == 16) begin
					state<=5;
					out<=244;
				end
				if(in == 17) begin
					state<=5;
					out<=245;
				end
				if(in == 18) begin
					state<=5;
					out<=246;
				end
				if(in == 19) begin
					state<=5;
					out<=247;
				end
				if(in == 20) begin
					state<=5;
					out<=248;
				end
				if(in == 21) begin
					state<=5;
					out<=249;
				end
				if(in == 22) begin
					state<=5;
					out<=250;
				end
				if(in == 23) begin
					state<=5;
					out<=251;
				end
				if(in == 24) begin
					state<=5;
					out<=252;
				end
				if(in == 25) begin
					state<=5;
					out<=253;
				end
				if(in == 26) begin
					state<=5;
					out<=254;
				end
				if(in == 27) begin
					state<=5;
					out<=255;
				end
				if(in == 28) begin
					state<=5;
					out<=0;
				end
				if(in == 29) begin
					state<=5;
					out<=1;
				end
				if(in == 30) begin
					state<=5;
					out<=2;
				end
				if(in == 31) begin
					state<=5;
					out<=3;
				end
				if(in == 32) begin
					state<=5;
					out<=4;
				end
				if(in == 33) begin
					state<=5;
					out<=5;
				end
				if(in == 34) begin
					state<=5;
					out<=6;
				end
				if(in == 35) begin
					state<=5;
					out<=7;
				end
				if(in == 36) begin
					state<=5;
					out<=8;
				end
				if(in == 37) begin
					state<=5;
					out<=9;
				end
				if(in == 38) begin
					state<=5;
					out<=10;
				end
				if(in == 39) begin
					state<=5;
					out<=11;
				end
				if(in == 40) begin
					state<=5;
					out<=12;
				end
				if(in == 41) begin
					state<=5;
					out<=13;
				end
				if(in == 42) begin
					state<=5;
					out<=14;
				end
				if(in == 43) begin
					state<=5;
					out<=15;
				end
				if(in == 44) begin
					state<=5;
					out<=16;
				end
				if(in == 45) begin
					state<=5;
					out<=17;
				end
				if(in == 46) begin
					state<=5;
					out<=18;
				end
				if(in == 47) begin
					state<=5;
					out<=19;
				end
				if(in == 48) begin
					state<=5;
					out<=20;
				end
				if(in == 49) begin
					state<=5;
					out<=21;
				end
				if(in == 50) begin
					state<=5;
					out<=22;
				end
				if(in == 51) begin
					state<=5;
					out<=23;
				end
				if(in == 52) begin
					state<=5;
					out<=24;
				end
				if(in == 53) begin
					state<=3;
					out<=25;
				end
				if(in == 54) begin
					state<=4;
					out<=26;
				end
				if(in == 55) begin
					state<=3;
					out<=27;
				end
				if(in == 56) begin
					state<=5;
					out<=28;
				end
				if(in == 57) begin
					state<=3;
					out<=29;
				end
				if(in == 58) begin
					state<=5;
					out<=30;
				end
				if(in == 59) begin
					state<=5;
					out<=31;
				end
				if(in == 60) begin
					state<=5;
					out<=32;
				end
				if(in == 61) begin
					state<=5;
					out<=33;
				end
				if(in == 62) begin
					state<=5;
					out<=34;
				end
				if(in == 63) begin
					state<=5;
					out<=35;
				end
				if(in == 64) begin
					state<=5;
					out<=36;
				end
				if(in == 65) begin
					state<=5;
					out<=37;
				end
				if(in == 66) begin
					state<=5;
					out<=38;
				end
				if(in == 67) begin
					state<=5;
					out<=39;
				end
				if(in == 68) begin
					state<=5;
					out<=40;
				end
				if(in == 69) begin
					state<=5;
					out<=41;
				end
				if(in == 70) begin
					state<=5;
					out<=42;
				end
				if(in == 71) begin
					state<=5;
					out<=43;
				end
				if(in == 72) begin
					state<=5;
					out<=44;
				end
				if(in == 73) begin
					state<=5;
					out<=45;
				end
				if(in == 74) begin
					state<=5;
					out<=46;
				end
				if(in == 75) begin
					state<=5;
					out<=47;
				end
				if(in == 76) begin
					state<=5;
					out<=48;
				end
				if(in == 77) begin
					state<=5;
					out<=49;
				end
				if(in == 78) begin
					state<=5;
					out<=50;
				end
				if(in == 79) begin
					state<=5;
					out<=51;
				end
				if(in == 80) begin
					state<=5;
					out<=52;
				end
				if(in == 81) begin
					state<=5;
					out<=53;
				end
				if(in == 82) begin
					state<=5;
					out<=54;
				end
				if(in == 83) begin
					state<=5;
					out<=55;
				end
				if(in == 84) begin
					state<=5;
					out<=56;
				end
				if(in == 85) begin
					state<=5;
					out<=57;
				end
				if(in == 86) begin
					state<=5;
					out<=58;
				end
				if(in == 87) begin
					state<=5;
					out<=59;
				end
				if(in == 88) begin
					state<=5;
					out<=60;
				end
				if(in == 89) begin
					state<=5;
					out<=61;
				end
				if(in == 90) begin
					state<=5;
					out<=62;
				end
				if(in == 91) begin
					state<=5;
					out<=63;
				end
				if(in == 92) begin
					state<=5;
					out<=64;
				end
				if(in == 93) begin
					state<=5;
					out<=65;
				end
				if(in == 94) begin
					state<=5;
					out<=66;
				end
				if(in == 95) begin
					state<=5;
					out<=67;
				end
				if(in == 96) begin
					state<=5;
					out<=68;
				end
				if(in == 97) begin
					state<=5;
					out<=69;
				end
				if(in == 98) begin
					state<=5;
					out<=70;
				end
				if(in == 99) begin
					state<=5;
					out<=71;
				end
				if(in == 100) begin
					state<=5;
					out<=72;
				end
				if(in == 101) begin
					state<=5;
					out<=73;
				end
				if(in == 102) begin
					state<=5;
					out<=74;
				end
				if(in == 103) begin
					state<=5;
					out<=75;
				end
				if(in == 104) begin
					state<=5;
					out<=76;
				end
				if(in == 105) begin
					state<=2;
					out<=77;
				end
				if(in == 106) begin
					state<=2;
					out<=78;
				end
				if(in == 107) begin
					state<=2;
					out<=79;
				end
				if(in == 108) begin
					state<=2;
					out<=80;
				end
				if(in == 109) begin
					state<=2;
					out<=81;
				end
				if(in == 110) begin
					state<=2;
					out<=82;
				end
				if(in == 111) begin
					state<=2;
					out<=83;
				end
				if(in == 112) begin
					state<=2;
					out<=84;
				end
				if(in == 113) begin
					state<=2;
					out<=85;
				end
				if(in == 114) begin
					state<=2;
					out<=86;
				end
				if(in == 115) begin
					state<=2;
					out<=87;
				end
				if(in == 116) begin
					state<=2;
					out<=88;
				end
				if(in == 117) begin
					state<=3;
					out<=89;
				end
				if(in == 118) begin
					state<=4;
					out<=90;
				end
				if(in == 119) begin
					state<=3;
					out<=91;
				end
				if(in == 120) begin
					state<=5;
					out<=92;
				end
				if(in == 121) begin
					state<=3;
					out<=93;
				end
				if(in == 122) begin
					state<=5;
					out<=94;
				end
				if(in == 123) begin
					state<=5;
					out<=95;
				end
				if(in == 124) begin
					state<=5;
					out<=96;
				end
				if(in == 125) begin
					state<=5;
					out<=97;
				end
				if(in == 126) begin
					state<=5;
					out<=98;
				end
				if(in == 127) begin
					state<=5;
					out<=99;
				end
				if(in == 128) begin
					state<=5;
					out<=100;
				end
				if(in == 129) begin
					state<=5;
					out<=101;
				end
				if(in == 130) begin
					state<=5;
					out<=102;
				end
				if(in == 131) begin
					state<=5;
					out<=103;
				end
				if(in == 132) begin
					state<=5;
					out<=104;
				end
				if(in == 133) begin
					state<=5;
					out<=105;
				end
				if(in == 134) begin
					state<=5;
					out<=106;
				end
				if(in == 135) begin
					state<=5;
					out<=107;
				end
				if(in == 136) begin
					state<=5;
					out<=108;
				end
				if(in == 137) begin
					state<=5;
					out<=109;
				end
				if(in == 138) begin
					state<=5;
					out<=110;
				end
				if(in == 139) begin
					state<=5;
					out<=111;
				end
				if(in == 140) begin
					state<=5;
					out<=112;
				end
				if(in == 141) begin
					state<=5;
					out<=113;
				end
				if(in == 142) begin
					state<=5;
					out<=114;
				end
				if(in == 143) begin
					state<=5;
					out<=115;
				end
				if(in == 144) begin
					state<=5;
					out<=116;
				end
				if(in == 145) begin
					state<=5;
					out<=117;
				end
				if(in == 146) begin
					state<=5;
					out<=118;
				end
				if(in == 147) begin
					state<=5;
					out<=119;
				end
				if(in == 148) begin
					state<=5;
					out<=120;
				end
				if(in == 149) begin
					state<=5;
					out<=121;
				end
				if(in == 150) begin
					state<=5;
					out<=122;
				end
				if(in == 151) begin
					state<=5;
					out<=123;
				end
				if(in == 152) begin
					state<=5;
					out<=124;
				end
				if(in == 153) begin
					state<=5;
					out<=125;
				end
				if(in == 154) begin
					state<=5;
					out<=126;
				end
				if(in == 155) begin
					state<=5;
					out<=127;
				end
				if(in == 156) begin
					state<=5;
					out<=128;
				end
				if(in == 157) begin
					state<=5;
					out<=129;
				end
				if(in == 158) begin
					state<=5;
					out<=130;
				end
				if(in == 159) begin
					state<=5;
					out<=131;
				end
				if(in == 160) begin
					state<=5;
					out<=132;
				end
				if(in == 161) begin
					state<=5;
					out<=133;
				end
				if(in == 162) begin
					state<=5;
					out<=134;
				end
				if(in == 163) begin
					state<=5;
					out<=135;
				end
				if(in == 164) begin
					state<=5;
					out<=136;
				end
				if(in == 165) begin
					state<=5;
					out<=137;
				end
				if(in == 166) begin
					state<=5;
					out<=138;
				end
				if(in == 167) begin
					state<=5;
					out<=139;
				end
				if(in == 168) begin
					state<=5;
					out<=140;
				end
				if(in == 169) begin
					state<=3;
					out<=141;
				end
				if(in == 170) begin
					state<=4;
					out<=142;
				end
				if(in == 171) begin
					state<=3;
					out<=143;
				end
				if(in == 172) begin
					state<=5;
					out<=144;
				end
				if(in == 173) begin
					state<=3;
					out<=145;
				end
				if(in == 174) begin
					state<=5;
					out<=146;
				end
				if(in == 175) begin
					state<=5;
					out<=147;
				end
				if(in == 176) begin
					state<=5;
					out<=148;
				end
				if(in == 177) begin
					state<=5;
					out<=149;
				end
				if(in == 178) begin
					state<=5;
					out<=150;
				end
				if(in == 179) begin
					state<=5;
					out<=151;
				end
				if(in == 180) begin
					state<=5;
					out<=152;
				end
				if(in == 181) begin
					state<=5;
					out<=153;
				end
				if(in == 182) begin
					state<=5;
					out<=154;
				end
				if(in == 183) begin
					state<=5;
					out<=155;
				end
				if(in == 184) begin
					state<=5;
					out<=156;
				end
				if(in == 185) begin
					state<=5;
					out<=157;
				end
				if(in == 186) begin
					state<=5;
					out<=158;
				end
				if(in == 187) begin
					state<=5;
					out<=159;
				end
				if(in == 188) begin
					state<=5;
					out<=160;
				end
				if(in == 189) begin
					state<=5;
					out<=161;
				end
				if(in == 190) begin
					state<=5;
					out<=162;
				end
				if(in == 191) begin
					state<=5;
					out<=163;
				end
				if(in == 192) begin
					state<=5;
					out<=164;
				end
				if(in == 193) begin
					state<=5;
					out<=165;
				end
				if(in == 194) begin
					state<=5;
					out<=166;
				end
				if(in == 195) begin
					state<=5;
					out<=167;
				end
				if(in == 196) begin
					state<=5;
					out<=168;
				end
				if(in == 197) begin
					state<=5;
					out<=169;
				end
				if(in == 198) begin
					state<=5;
					out<=170;
				end
				if(in == 199) begin
					state<=5;
					out<=171;
				end
				if(in == 200) begin
					state<=5;
					out<=172;
				end
				if(in == 201) begin
					state<=5;
					out<=173;
				end
				if(in == 202) begin
					state<=5;
					out<=174;
				end
				if(in == 203) begin
					state<=5;
					out<=175;
				end
				if(in == 204) begin
					state<=5;
					out<=176;
				end
				if(in == 205) begin
					state<=5;
					out<=177;
				end
				if(in == 206) begin
					state<=5;
					out<=178;
				end
				if(in == 207) begin
					state<=5;
					out<=179;
				end
				if(in == 208) begin
					state<=5;
					out<=180;
				end
				if(in == 209) begin
					state<=5;
					out<=181;
				end
				if(in == 210) begin
					state<=5;
					out<=182;
				end
				if(in == 211) begin
					state<=5;
					out<=183;
				end
				if(in == 212) begin
					state<=5;
					out<=184;
				end
				if(in == 213) begin
					state<=5;
					out<=185;
				end
				if(in == 214) begin
					state<=5;
					out<=186;
				end
				if(in == 215) begin
					state<=5;
					out<=187;
				end
				if(in == 216) begin
					state<=5;
					out<=188;
				end
				if(in == 217) begin
					state<=5;
					out<=189;
				end
				if(in == 218) begin
					state<=5;
					out<=190;
				end
				if(in == 219) begin
					state<=5;
					out<=191;
				end
				if(in == 220) begin
					state<=5;
					out<=192;
				end
				if(in == 221) begin
					state<=2;
					out<=193;
				end
				if(in == 222) begin
					state<=2;
					out<=194;
				end
				if(in == 223) begin
					state<=2;
					out<=195;
				end
				if(in == 224) begin
					state<=2;
					out<=196;
				end
				if(in == 225) begin
					state<=2;
					out<=197;
				end
				if(in == 226) begin
					state<=2;
					out<=198;
				end
				if(in == 227) begin
					state<=2;
					out<=199;
				end
				if(in == 228) begin
					state<=2;
					out<=200;
				end
				if(in == 229) begin
					state<=2;
					out<=201;
				end
				if(in == 230) begin
					state<=2;
					out<=202;
				end
				if(in == 231) begin
					state<=2;
					out<=203;
				end
				if(in == 232) begin
					state<=2;
					out<=204;
				end
				if(in == 233) begin
					state<=3;
					out<=205;
				end
				if(in == 234) begin
					state<=4;
					out<=206;
				end
				if(in == 235) begin
					state<=3;
					out<=207;
				end
				if(in == 236) begin
					state<=5;
					out<=208;
				end
				if(in == 237) begin
					state<=3;
					out<=209;
				end
				if(in == 238) begin
					state<=5;
					out<=210;
				end
				if(in == 239) begin
					state<=5;
					out<=211;
				end
				if(in == 240) begin
					state<=5;
					out<=212;
				end
				if(in == 241) begin
					state<=5;
					out<=213;
				end
				if(in == 242) begin
					state<=5;
					out<=214;
				end
				if(in == 243) begin
					state<=5;
					out<=215;
				end
				if(in == 244) begin
					state<=5;
					out<=216;
				end
				if(in == 245) begin
					state<=5;
					out<=217;
				end
				if(in == 246) begin
					state<=5;
					out<=218;
				end
				if(in == 247) begin
					state<=5;
					out<=219;
				end
				if(in == 248) begin
					state<=5;
					out<=220;
				end
				if(in == 249) begin
					state<=5;
					out<=221;
				end
				if(in == 250) begin
					state<=5;
					out<=222;
				end
				if(in == 251) begin
					state<=5;
					out<=223;
				end
				if(in == 252) begin
					state<=5;
					out<=224;
				end
				if(in == 253) begin
					state<=5;
					out<=225;
				end
				if(in == 254) begin
					state<=5;
					out<=226;
				end
				if(in == 255) begin
					state<=5;
					out<=227;
				end
				if(in == 256) begin
					state<=5;
					out<=228;
				end
				if(in == 257) begin
					state<=5;
					out<=229;
				end
				if(in == 258) begin
					state<=5;
					out<=230;
				end
				if(in == 259) begin
					state<=5;
					out<=231;
				end
				if(in == 260) begin
					state<=5;
					out<=232;
				end
				if(in == 261) begin
					state<=5;
					out<=233;
				end
				if(in == 262) begin
					state<=5;
					out<=234;
				end
				if(in == 263) begin
					state<=5;
					out<=235;
				end
				if(in == 264) begin
					state<=5;
					out<=236;
				end
				if(in == 265) begin
					state<=5;
					out<=237;
				end
				if(in == 266) begin
					state<=5;
					out<=238;
				end
				if(in == 267) begin
					state<=5;
					out<=239;
				end
				if(in == 268) begin
					state<=5;
					out<=240;
				end
				if(in == 269) begin
					state<=5;
					out<=241;
				end
				if(in == 270) begin
					state<=5;
					out<=242;
				end
				if(in == 271) begin
					state<=5;
					out<=243;
				end
				if(in == 272) begin
					state<=5;
					out<=244;
				end
				if(in == 273) begin
					state<=5;
					out<=245;
				end
				if(in == 274) begin
					state<=5;
					out<=246;
				end
				if(in == 275) begin
					state<=5;
					out<=247;
				end
				if(in == 276) begin
					state<=5;
					out<=248;
				end
				if(in == 277) begin
					state<=5;
					out<=249;
				end
				if(in == 278) begin
					state<=5;
					out<=250;
				end
				if(in == 279) begin
					state<=5;
					out<=251;
				end
				if(in == 280) begin
					state<=5;
					out<=252;
				end
				if(in == 281) begin
					state<=5;
					out<=253;
				end
				if(in == 282) begin
					state<=5;
					out<=254;
				end
				if(in == 283) begin
					state<=5;
					out<=255;
				end
				if(in == 284) begin
					state<=5;
					out<=0;
				end
				if(in == 285) begin
					state<=3;
					out<=1;
				end
				if(in == 286) begin
					state<=4;
					out<=2;
				end
				if(in == 287) begin
					state<=3;
					out<=3;
				end
				if(in == 288) begin
					state<=5;
					out<=4;
				end
				if(in == 289) begin
					state<=3;
					out<=5;
				end
				if(in == 290) begin
					state<=5;
					out<=6;
				end
				if(in == 291) begin
					state<=5;
					out<=7;
				end
				if(in == 292) begin
					state<=5;
					out<=8;
				end
				if(in == 293) begin
					state<=5;
					out<=9;
				end
				if(in == 294) begin
					state<=5;
					out<=10;
				end
				if(in == 295) begin
					state<=5;
					out<=11;
				end
				if(in == 296) begin
					state<=5;
					out<=12;
				end
				if(in == 297) begin
					state<=5;
					out<=13;
				end
				if(in == 298) begin
					state<=5;
					out<=14;
				end
				if(in == 299) begin
					state<=5;
					out<=15;
				end
				if(in == 300) begin
					state<=5;
					out<=16;
				end
				if(in == 301) begin
					state<=5;
					out<=17;
				end
				if(in == 302) begin
					state<=5;
					out<=18;
				end
				if(in == 303) begin
					state<=5;
					out<=19;
				end
				if(in == 304) begin
					state<=5;
					out<=20;
				end
				if(in == 305) begin
					state<=5;
					out<=21;
				end
				if(in == 306) begin
					state<=5;
					out<=22;
				end
				if(in == 307) begin
					state<=5;
					out<=23;
				end
				if(in == 308) begin
					state<=5;
					out<=24;
				end
				if(in == 309) begin
					state<=5;
					out<=25;
				end
				if(in == 310) begin
					state<=5;
					out<=26;
				end
				if(in == 311) begin
					state<=5;
					out<=27;
				end
				if(in == 312) begin
					state<=5;
					out<=28;
				end
				if(in == 313) begin
					state<=5;
					out<=29;
				end
				if(in == 314) begin
					state<=5;
					out<=30;
				end
				if(in == 315) begin
					state<=5;
					out<=31;
				end
				if(in == 316) begin
					state<=5;
					out<=32;
				end
				if(in == 317) begin
					state<=5;
					out<=33;
				end
				if(in == 318) begin
					state<=5;
					out<=34;
				end
				if(in == 319) begin
					state<=5;
					out<=35;
				end
				if(in == 320) begin
					state<=5;
					out<=36;
				end
				if(in == 321) begin
					state<=5;
					out<=37;
				end
				if(in == 322) begin
					state<=5;
					out<=38;
				end
				if(in == 323) begin
					state<=5;
					out<=39;
				end
				if(in == 324) begin
					state<=5;
					out<=40;
				end
				if(in == 325) begin
					state<=5;
					out<=41;
				end
				if(in == 326) begin
					state<=5;
					out<=42;
				end
				if(in == 327) begin
					state<=5;
					out<=43;
				end
				if(in == 328) begin
					state<=5;
					out<=44;
				end
				if(in == 329) begin
					state<=5;
					out<=45;
				end
				if(in == 330) begin
					state<=5;
					out<=46;
				end
				if(in == 331) begin
					state<=5;
					out<=47;
				end
				if(in == 332) begin
					state<=5;
					out<=48;
				end
				if(in == 333) begin
					state<=5;
					out<=49;
				end
				if(in == 334) begin
					state<=5;
					out<=50;
				end
				if(in == 335) begin
					state<=5;
					out<=51;
				end
				if(in == 336) begin
					state<=5;
					out<=52;
				end
				if(in == 337) begin
					state<=2;
					out<=53;
				end
				if(in == 338) begin
					state<=2;
					out<=54;
				end
				if(in == 339) begin
					state<=2;
					out<=55;
				end
				if(in == 340) begin
					state<=2;
					out<=56;
				end
				if(in == 341) begin
					state<=2;
					out<=57;
				end
				if(in == 342) begin
					state<=2;
					out<=58;
				end
				if(in == 343) begin
					state<=2;
					out<=59;
				end
				if(in == 344) begin
					state<=2;
					out<=60;
				end
				if(in == 345) begin
					state<=2;
					out<=61;
				end
				if(in == 346) begin
					state<=2;
					out<=62;
				end
				if(in == 347) begin
					state<=2;
					out<=63;
				end
				if(in == 348) begin
					state<=2;
					out<=64;
				end
				if(in == 349) begin
					state<=3;
					out<=65;
				end
				if(in == 350) begin
					state<=4;
					out<=66;
				end
				if(in == 351) begin
					state<=3;
					out<=67;
				end
				if(in == 352) begin
					state<=5;
					out<=68;
				end
				if(in == 353) begin
					state<=3;
					out<=69;
				end
				if(in == 354) begin
					state<=5;
					out<=70;
				end
				if(in == 355) begin
					state<=5;
					out<=71;
				end
				if(in == 356) begin
					state<=5;
					out<=72;
				end
				if(in == 357) begin
					state<=5;
					out<=73;
				end
				if(in == 358) begin
					state<=5;
					out<=74;
				end
				if(in == 359) begin
					state<=5;
					out<=75;
				end
				if(in == 360) begin
					state<=5;
					out<=76;
				end
				if(in == 361) begin
					state<=5;
					out<=77;
				end
				if(in == 362) begin
					state<=5;
					out<=78;
				end
				if(in == 363) begin
					state<=5;
					out<=79;
				end
				if(in == 364) begin
					state<=5;
					out<=80;
				end
				if(in == 365) begin
					state<=5;
					out<=81;
				end
				if(in == 366) begin
					state<=5;
					out<=82;
				end
				if(in == 367) begin
					state<=5;
					out<=83;
				end
				if(in == 368) begin
					state<=5;
					out<=84;
				end
				if(in == 369) begin
					state<=5;
					out<=85;
				end
				if(in == 370) begin
					state<=5;
					out<=86;
				end
				if(in == 371) begin
					state<=5;
					out<=87;
				end
				if(in == 372) begin
					state<=5;
					out<=88;
				end
				if(in == 373) begin
					state<=5;
					out<=89;
				end
				if(in == 374) begin
					state<=5;
					out<=90;
				end
				if(in == 375) begin
					state<=5;
					out<=91;
				end
				if(in == 376) begin
					state<=5;
					out<=92;
				end
				if(in == 377) begin
					state<=5;
					out<=93;
				end
				if(in == 378) begin
					state<=5;
					out<=94;
				end
				if(in == 379) begin
					state<=5;
					out<=95;
				end
				if(in == 380) begin
					state<=5;
					out<=96;
				end
				if(in == 381) begin
					state<=5;
					out<=97;
				end
				if(in == 382) begin
					state<=5;
					out<=98;
				end
				if(in == 383) begin
					state<=5;
					out<=99;
				end
				if(in == 384) begin
					state<=5;
					out<=100;
				end
				if(in == 385) begin
					state<=5;
					out<=101;
				end
				if(in == 386) begin
					state<=5;
					out<=102;
				end
				if(in == 387) begin
					state<=5;
					out<=103;
				end
				if(in == 388) begin
					state<=5;
					out<=104;
				end
				if(in == 389) begin
					state<=5;
					out<=105;
				end
				if(in == 390) begin
					state<=5;
					out<=106;
				end
				if(in == 391) begin
					state<=5;
					out<=107;
				end
				if(in == 392) begin
					state<=5;
					out<=108;
				end
				if(in == 393) begin
					state<=5;
					out<=109;
				end
				if(in == 394) begin
					state<=5;
					out<=110;
				end
				if(in == 395) begin
					state<=5;
					out<=111;
				end
				if(in == 396) begin
					state<=5;
					out<=112;
				end
				if(in == 397) begin
					state<=5;
					out<=113;
				end
				if(in == 398) begin
					state<=5;
					out<=114;
				end
				if(in == 399) begin
					state<=5;
					out<=115;
				end
				if(in == 400) begin
					state<=5;
					out<=116;
				end
				if(in == 401) begin
					state<=3;
					out<=117;
				end
				if(in == 402) begin
					state<=4;
					out<=118;
				end
				if(in == 403) begin
					state<=3;
					out<=119;
				end
				if(in == 404) begin
					state<=5;
					out<=120;
				end
				if(in == 405) begin
					state<=3;
					out<=121;
				end
				if(in == 406) begin
					state<=5;
					out<=122;
				end
				if(in == 407) begin
					state<=5;
					out<=123;
				end
				if(in == 408) begin
					state<=5;
					out<=124;
				end
				if(in == 409) begin
					state<=5;
					out<=125;
				end
				if(in == 410) begin
					state<=5;
					out<=126;
				end
				if(in == 411) begin
					state<=5;
					out<=127;
				end
				if(in == 412) begin
					state<=5;
					out<=128;
				end
				if(in == 413) begin
					state<=5;
					out<=129;
				end
				if(in == 414) begin
					state<=5;
					out<=130;
				end
				if(in == 415) begin
					state<=5;
					out<=131;
				end
				if(in == 416) begin
					state<=5;
					out<=132;
				end
				if(in == 417) begin
					state<=5;
					out<=133;
				end
				if(in == 418) begin
					state<=5;
					out<=134;
				end
				if(in == 419) begin
					state<=5;
					out<=135;
				end
				if(in == 420) begin
					state<=5;
					out<=136;
				end
				if(in == 421) begin
					state<=5;
					out<=137;
				end
				if(in == 422) begin
					state<=5;
					out<=138;
				end
				if(in == 423) begin
					state<=5;
					out<=139;
				end
				if(in == 424) begin
					state<=5;
					out<=140;
				end
				if(in == 425) begin
					state<=5;
					out<=141;
				end
				if(in == 426) begin
					state<=5;
					out<=142;
				end
				if(in == 427) begin
					state<=5;
					out<=143;
				end
				if(in == 428) begin
					state<=5;
					out<=144;
				end
				if(in == 429) begin
					state<=5;
					out<=145;
				end
				if(in == 430) begin
					state<=5;
					out<=146;
				end
				if(in == 431) begin
					state<=5;
					out<=147;
				end
				if(in == 432) begin
					state<=5;
					out<=148;
				end
				if(in == 433) begin
					state<=5;
					out<=149;
				end
				if(in == 434) begin
					state<=5;
					out<=150;
				end
				if(in == 435) begin
					state<=5;
					out<=151;
				end
				if(in == 436) begin
					state<=5;
					out<=152;
				end
				if(in == 437) begin
					state<=5;
					out<=153;
				end
				if(in == 438) begin
					state<=5;
					out<=154;
				end
				if(in == 439) begin
					state<=5;
					out<=155;
				end
				if(in == 440) begin
					state<=5;
					out<=156;
				end
				if(in == 441) begin
					state<=5;
					out<=157;
				end
				if(in == 442) begin
					state<=5;
					out<=158;
				end
				if(in == 443) begin
					state<=5;
					out<=159;
				end
				if(in == 444) begin
					state<=5;
					out<=160;
				end
				if(in == 445) begin
					state<=5;
					out<=161;
				end
				if(in == 446) begin
					state<=5;
					out<=162;
				end
				if(in == 447) begin
					state<=5;
					out<=163;
				end
				if(in == 448) begin
					state<=5;
					out<=164;
				end
				if(in == 449) begin
					state<=5;
					out<=165;
				end
				if(in == 450) begin
					state<=5;
					out<=166;
				end
				if(in == 451) begin
					state<=5;
					out<=167;
				end
				if(in == 452) begin
					state<=5;
					out<=168;
				end
				if(in == 453) begin
					state<=2;
					out<=169;
				end
				if(in == 454) begin
					state<=2;
					out<=170;
				end
				if(in == 455) begin
					state<=2;
					out<=171;
				end
				if(in == 456) begin
					state<=2;
					out<=172;
				end
				if(in == 457) begin
					state<=2;
					out<=173;
				end
				if(in == 458) begin
					state<=2;
					out<=174;
				end
				if(in == 459) begin
					state<=2;
					out<=175;
				end
				if(in == 460) begin
					state<=2;
					out<=176;
				end
				if(in == 461) begin
					state<=2;
					out<=177;
				end
				if(in == 462) begin
					state<=2;
					out<=178;
				end
				if(in == 463) begin
					state<=2;
					out<=179;
				end
				if(in == 464) begin
					state<=2;
					out<=180;
				end
				if(in == 465) begin
					state<=3;
					out<=181;
				end
				if(in == 466) begin
					state<=4;
					out<=182;
				end
				if(in == 467) begin
					state<=3;
					out<=183;
				end
				if(in == 468) begin
					state<=5;
					out<=184;
				end
				if(in == 469) begin
					state<=3;
					out<=185;
				end
				if(in == 470) begin
					state<=5;
					out<=186;
				end
				if(in == 471) begin
					state<=5;
					out<=187;
				end
				if(in == 472) begin
					state<=5;
					out<=188;
				end
				if(in == 473) begin
					state<=5;
					out<=189;
				end
				if(in == 474) begin
					state<=5;
					out<=190;
				end
				if(in == 475) begin
					state<=5;
					out<=191;
				end
				if(in == 476) begin
					state<=5;
					out<=192;
				end
				if(in == 477) begin
					state<=5;
					out<=193;
				end
				if(in == 478) begin
					state<=5;
					out<=194;
				end
				if(in == 479) begin
					state<=5;
					out<=195;
				end
				if(in == 480) begin
					state<=5;
					out<=196;
				end
				if(in == 481) begin
					state<=5;
					out<=197;
				end
				if(in == 482) begin
					state<=5;
					out<=198;
				end
				if(in == 483) begin
					state<=5;
					out<=199;
				end
				if(in == 484) begin
					state<=5;
					out<=200;
				end
				if(in == 485) begin
					state<=5;
					out<=201;
				end
				if(in == 486) begin
					state<=5;
					out<=202;
				end
				if(in == 487) begin
					state<=5;
					out<=203;
				end
				if(in == 488) begin
					state<=5;
					out<=204;
				end
				if(in == 489) begin
					state<=5;
					out<=205;
				end
				if(in == 490) begin
					state<=5;
					out<=206;
				end
				if(in == 491) begin
					state<=5;
					out<=207;
				end
				if(in == 492) begin
					state<=5;
					out<=208;
				end
				if(in == 493) begin
					state<=5;
					out<=209;
				end
				if(in == 494) begin
					state<=5;
					out<=210;
				end
				if(in == 495) begin
					state<=5;
					out<=211;
				end
				if(in == 496) begin
					state<=5;
					out<=212;
				end
				if(in == 497) begin
					state<=5;
					out<=213;
				end
				if(in == 498) begin
					state<=5;
					out<=214;
				end
				if(in == 499) begin
					state<=5;
					out<=215;
				end
				if(in == 500) begin
					state<=5;
					out<=216;
				end
				if(in == 501) begin
					state<=5;
					out<=217;
				end
				if(in == 502) begin
					state<=5;
					out<=218;
				end
				if(in == 503) begin
					state<=5;
					out<=219;
				end
				if(in == 504) begin
					state<=5;
					out<=220;
				end
				if(in == 505) begin
					state<=5;
					out<=221;
				end
				if(in == 506) begin
					state<=5;
					out<=222;
				end
				if(in == 507) begin
					state<=5;
					out<=223;
				end
				if(in == 508) begin
					state<=5;
					out<=224;
				end
				if(in == 509) begin
					state<=5;
					out<=225;
				end
				if(in == 510) begin
					state<=5;
					out<=226;
				end
				if(in == 511) begin
					state<=5;
					out<=227;
				end
				if(in == 512) begin
					state<=5;
					out<=228;
				end
				if(in == 513) begin
					state<=5;
					out<=229;
				end
				if(in == 514) begin
					state<=5;
					out<=230;
				end
				if(in == 515) begin
					state<=5;
					out<=231;
				end
				if(in == 516) begin
					state<=5;
					out<=232;
				end
				if(in == 517) begin
					state<=3;
					out<=233;
				end
				if(in == 518) begin
					state<=4;
					out<=234;
				end
				if(in == 519) begin
					state<=3;
					out<=235;
				end
				if(in == 520) begin
					state<=5;
					out<=236;
				end
				if(in == 521) begin
					state<=3;
					out<=237;
				end
				if(in == 522) begin
					state<=5;
					out<=238;
				end
				if(in == 523) begin
					state<=5;
					out<=239;
				end
				if(in == 524) begin
					state<=5;
					out<=240;
				end
				if(in == 525) begin
					state<=5;
					out<=241;
				end
				if(in == 526) begin
					state<=5;
					out<=242;
				end
				if(in == 527) begin
					state<=5;
					out<=243;
				end
				if(in == 528) begin
					state<=5;
					out<=244;
				end
				if(in == 529) begin
					state<=5;
					out<=245;
				end
				if(in == 530) begin
					state<=5;
					out<=246;
				end
				if(in == 531) begin
					state<=5;
					out<=247;
				end
				if(in == 532) begin
					state<=5;
					out<=248;
				end
				if(in == 533) begin
					state<=5;
					out<=249;
				end
				if(in == 534) begin
					state<=5;
					out<=250;
				end
				if(in == 535) begin
					state<=5;
					out<=251;
				end
				if(in == 536) begin
					state<=5;
					out<=252;
				end
				if(in == 537) begin
					state<=5;
					out<=253;
				end
				if(in == 538) begin
					state<=5;
					out<=254;
				end
				if(in == 539) begin
					state<=5;
					out<=255;
				end
				if(in == 540) begin
					state<=5;
					out<=0;
				end
				if(in == 541) begin
					state<=5;
					out<=1;
				end
				if(in == 542) begin
					state<=5;
					out<=2;
				end
				if(in == 543) begin
					state<=5;
					out<=3;
				end
				if(in == 544) begin
					state<=5;
					out<=4;
				end
				if(in == 545) begin
					state<=5;
					out<=5;
				end
				if(in == 546) begin
					state<=5;
					out<=6;
				end
				if(in == 547) begin
					state<=5;
					out<=7;
				end
				if(in == 548) begin
					state<=5;
					out<=8;
				end
				if(in == 549) begin
					state<=5;
					out<=9;
				end
				if(in == 550) begin
					state<=5;
					out<=10;
				end
				if(in == 551) begin
					state<=5;
					out<=11;
				end
				if(in == 552) begin
					state<=5;
					out<=12;
				end
				if(in == 553) begin
					state<=5;
					out<=13;
				end
				if(in == 554) begin
					state<=5;
					out<=14;
				end
				if(in == 555) begin
					state<=5;
					out<=15;
				end
				if(in == 556) begin
					state<=5;
					out<=16;
				end
				if(in == 557) begin
					state<=5;
					out<=17;
				end
				if(in == 558) begin
					state<=5;
					out<=18;
				end
				if(in == 559) begin
					state<=5;
					out<=19;
				end
				if(in == 560) begin
					state<=5;
					out<=20;
				end
				if(in == 561) begin
					state<=5;
					out<=21;
				end
				if(in == 562) begin
					state<=5;
					out<=22;
				end
				if(in == 563) begin
					state<=5;
					out<=23;
				end
				if(in == 564) begin
					state<=5;
					out<=24;
				end
				if(in == 565) begin
					state<=5;
					out<=25;
				end
				if(in == 566) begin
					state<=5;
					out<=26;
				end
				if(in == 567) begin
					state<=5;
					out<=27;
				end
				if(in == 568) begin
					state<=5;
					out<=28;
				end
				if(in == 569) begin
					state<=2;
					out<=29;
				end
				if(in == 570) begin
					state<=2;
					out<=30;
				end
				if(in == 571) begin
					state<=2;
					out<=31;
				end
				if(in == 572) begin
					state<=2;
					out<=32;
				end
				if(in == 573) begin
					state<=2;
					out<=33;
				end
				if(in == 574) begin
					state<=2;
					out<=34;
				end
				if(in == 575) begin
					state<=2;
					out<=35;
				end
				if(in == 576) begin
					state<=2;
					out<=36;
				end
				if(in == 577) begin
					state<=2;
					out<=37;
				end
				if(in == 578) begin
					state<=2;
					out<=38;
				end
				if(in == 579) begin
					state<=2;
					out<=39;
				end
				if(in == 580) begin
					state<=2;
					out<=40;
				end
				if(in == 581) begin
					state<=3;
					out<=41;
				end
				if(in == 582) begin
					state<=4;
					out<=42;
				end
				if(in == 583) begin
					state<=3;
					out<=43;
				end
				if(in == 584) begin
					state<=5;
					out<=44;
				end
				if(in == 585) begin
					state<=3;
					out<=45;
				end
				if(in == 586) begin
					state<=5;
					out<=46;
				end
				if(in == 587) begin
					state<=5;
					out<=47;
				end
				if(in == 588) begin
					state<=5;
					out<=48;
				end
				if(in == 589) begin
					state<=5;
					out<=49;
				end
				if(in == 590) begin
					state<=5;
					out<=50;
				end
				if(in == 591) begin
					state<=5;
					out<=51;
				end
				if(in == 592) begin
					state<=5;
					out<=52;
				end
				if(in == 593) begin
					state<=5;
					out<=53;
				end
				if(in == 594) begin
					state<=5;
					out<=54;
				end
				if(in == 595) begin
					state<=5;
					out<=55;
				end
				if(in == 596) begin
					state<=5;
					out<=56;
				end
				if(in == 597) begin
					state<=5;
					out<=57;
				end
				if(in == 598) begin
					state<=5;
					out<=58;
				end
				if(in == 599) begin
					state<=5;
					out<=59;
				end
				if(in == 600) begin
					state<=5;
					out<=60;
				end
				if(in == 601) begin
					state<=5;
					out<=61;
				end
				if(in == 602) begin
					state<=5;
					out<=62;
				end
				if(in == 603) begin
					state<=5;
					out<=63;
				end
				if(in == 604) begin
					state<=5;
					out<=64;
				end
				if(in == 605) begin
					state<=5;
					out<=65;
				end
				if(in == 606) begin
					state<=5;
					out<=66;
				end
				if(in == 607) begin
					state<=5;
					out<=67;
				end
				if(in == 608) begin
					state<=5;
					out<=68;
				end
				if(in == 609) begin
					state<=5;
					out<=69;
				end
				if(in == 610) begin
					state<=5;
					out<=70;
				end
				if(in == 611) begin
					state<=5;
					out<=71;
				end
				if(in == 612) begin
					state<=5;
					out<=72;
				end
				if(in == 613) begin
					state<=5;
					out<=73;
				end
				if(in == 614) begin
					state<=5;
					out<=74;
				end
				if(in == 615) begin
					state<=5;
					out<=75;
				end
				if(in == 616) begin
					state<=5;
					out<=76;
				end
				if(in == 617) begin
					state<=5;
					out<=77;
				end
				if(in == 618) begin
					state<=5;
					out<=78;
				end
				if(in == 619) begin
					state<=5;
					out<=79;
				end
				if(in == 620) begin
					state<=5;
					out<=80;
				end
				if(in == 621) begin
					state<=5;
					out<=81;
				end
				if(in == 622) begin
					state<=5;
					out<=82;
				end
				if(in == 623) begin
					state<=5;
					out<=83;
				end
				if(in == 624) begin
					state<=5;
					out<=84;
				end
				if(in == 625) begin
					state<=5;
					out<=85;
				end
				if(in == 626) begin
					state<=5;
					out<=86;
				end
				if(in == 627) begin
					state<=5;
					out<=87;
				end
				if(in == 628) begin
					state<=5;
					out<=88;
				end
				if(in == 629) begin
					state<=5;
					out<=89;
				end
				if(in == 630) begin
					state<=5;
					out<=90;
				end
				if(in == 631) begin
					state<=5;
					out<=91;
				end
				if(in == 632) begin
					state<=5;
					out<=92;
				end
				if(in == 633) begin
					state<=3;
					out<=93;
				end
				if(in == 634) begin
					state<=4;
					out<=94;
				end
				if(in == 635) begin
					state<=3;
					out<=95;
				end
				if(in == 636) begin
					state<=5;
					out<=96;
				end
				if(in == 637) begin
					state<=3;
					out<=97;
				end
				if(in == 638) begin
					state<=5;
					out<=98;
				end
				if(in == 639) begin
					state<=5;
					out<=99;
				end
				if(in == 640) begin
					state<=5;
					out<=100;
				end
				if(in == 641) begin
					state<=5;
					out<=101;
				end
				if(in == 642) begin
					state<=5;
					out<=102;
				end
				if(in == 643) begin
					state<=5;
					out<=103;
				end
				if(in == 644) begin
					state<=5;
					out<=104;
				end
				if(in == 645) begin
					state<=5;
					out<=105;
				end
				if(in == 646) begin
					state<=5;
					out<=106;
				end
				if(in == 647) begin
					state<=5;
					out<=107;
				end
				if(in == 648) begin
					state<=5;
					out<=108;
				end
				if(in == 649) begin
					state<=5;
					out<=109;
				end
				if(in == 650) begin
					state<=5;
					out<=110;
				end
				if(in == 651) begin
					state<=5;
					out<=111;
				end
				if(in == 652) begin
					state<=5;
					out<=112;
				end
				if(in == 653) begin
					state<=5;
					out<=113;
				end
				if(in == 654) begin
					state<=5;
					out<=114;
				end
				if(in == 655) begin
					state<=5;
					out<=115;
				end
				if(in == 656) begin
					state<=5;
					out<=116;
				end
				if(in == 657) begin
					state<=5;
					out<=117;
				end
				if(in == 658) begin
					state<=5;
					out<=118;
				end
				if(in == 659) begin
					state<=5;
					out<=119;
				end
				if(in == 660) begin
					state<=5;
					out<=120;
				end
				if(in == 661) begin
					state<=5;
					out<=121;
				end
				if(in == 662) begin
					state<=5;
					out<=122;
				end
				if(in == 663) begin
					state<=5;
					out<=123;
				end
				if(in == 664) begin
					state<=5;
					out<=124;
				end
				if(in == 665) begin
					state<=5;
					out<=125;
				end
				if(in == 666) begin
					state<=5;
					out<=126;
				end
				if(in == 667) begin
					state<=5;
					out<=127;
				end
				if(in == 668) begin
					state<=5;
					out<=128;
				end
				if(in == 669) begin
					state<=5;
					out<=129;
				end
				if(in == 670) begin
					state<=5;
					out<=130;
				end
				if(in == 671) begin
					state<=5;
					out<=131;
				end
				if(in == 672) begin
					state<=5;
					out<=132;
				end
				if(in == 673) begin
					state<=5;
					out<=133;
				end
				if(in == 674) begin
					state<=5;
					out<=134;
				end
				if(in == 675) begin
					state<=5;
					out<=135;
				end
				if(in == 676) begin
					state<=5;
					out<=136;
				end
				if(in == 677) begin
					state<=5;
					out<=137;
				end
				if(in == 678) begin
					state<=5;
					out<=138;
				end
				if(in == 679) begin
					state<=5;
					out<=139;
				end
				if(in == 680) begin
					state<=5;
					out<=140;
				end
				if(in == 681) begin
					state<=5;
					out<=141;
				end
				if(in == 682) begin
					state<=5;
					out<=142;
				end
				if(in == 683) begin
					state<=5;
					out<=143;
				end
				if(in == 684) begin
					state<=5;
					out<=144;
				end
				if(in == 685) begin
					state<=2;
					out<=145;
				end
				if(in == 686) begin
					state<=2;
					out<=146;
				end
				if(in == 687) begin
					state<=2;
					out<=147;
				end
				if(in == 688) begin
					state<=2;
					out<=148;
				end
				if(in == 689) begin
					state<=2;
					out<=149;
				end
				if(in == 690) begin
					state<=2;
					out<=150;
				end
				if(in == 691) begin
					state<=2;
					out<=151;
				end
				if(in == 692) begin
					state<=2;
					out<=152;
				end
				if(in == 693) begin
					state<=2;
					out<=153;
				end
				if(in == 694) begin
					state<=2;
					out<=154;
				end
				if(in == 695) begin
					state<=2;
					out<=155;
				end
				if(in == 696) begin
					state<=2;
					out<=156;
				end
				if(in == 697) begin
					state<=3;
					out<=157;
				end
				if(in == 698) begin
					state<=4;
					out<=158;
				end
				if(in == 699) begin
					state<=3;
					out<=159;
				end
				if(in == 700) begin
					state<=5;
					out<=160;
				end
				if(in == 701) begin
					state<=3;
					out<=161;
				end
				if(in == 702) begin
					state<=5;
					out<=162;
				end
				if(in == 703) begin
					state<=5;
					out<=163;
				end
				if(in == 704) begin
					state<=5;
					out<=164;
				end
				if(in == 705) begin
					state<=5;
					out<=165;
				end
				if(in == 706) begin
					state<=5;
					out<=166;
				end
				if(in == 707) begin
					state<=5;
					out<=167;
				end
				if(in == 708) begin
					state<=5;
					out<=168;
				end
				if(in == 709) begin
					state<=5;
					out<=169;
				end
				if(in == 710) begin
					state<=5;
					out<=170;
				end
				if(in == 711) begin
					state<=5;
					out<=171;
				end
				if(in == 712) begin
					state<=5;
					out<=172;
				end
				if(in == 713) begin
					state<=5;
					out<=173;
				end
				if(in == 714) begin
					state<=5;
					out<=174;
				end
				if(in == 715) begin
					state<=5;
					out<=175;
				end
				if(in == 716) begin
					state<=5;
					out<=176;
				end
				if(in == 717) begin
					state<=5;
					out<=177;
				end
				if(in == 718) begin
					state<=5;
					out<=178;
				end
				if(in == 719) begin
					state<=5;
					out<=179;
				end
				if(in == 720) begin
					state<=5;
					out<=180;
				end
				if(in == 721) begin
					state<=5;
					out<=181;
				end
				if(in == 722) begin
					state<=5;
					out<=182;
				end
				if(in == 723) begin
					state<=5;
					out<=183;
				end
				if(in == 724) begin
					state<=5;
					out<=184;
				end
				if(in == 725) begin
					state<=5;
					out<=185;
				end
				if(in == 726) begin
					state<=5;
					out<=186;
				end
				if(in == 727) begin
					state<=5;
					out<=187;
				end
				if(in == 728) begin
					state<=5;
					out<=188;
				end
				if(in == 729) begin
					state<=5;
					out<=189;
				end
				if(in == 730) begin
					state<=5;
					out<=190;
				end
				if(in == 731) begin
					state<=5;
					out<=191;
				end
				if(in == 732) begin
					state<=5;
					out<=192;
				end
				if(in == 733) begin
					state<=5;
					out<=193;
				end
				if(in == 734) begin
					state<=5;
					out<=194;
				end
				if(in == 735) begin
					state<=5;
					out<=195;
				end
				if(in == 736) begin
					state<=5;
					out<=196;
				end
				if(in == 737) begin
					state<=5;
					out<=197;
				end
				if(in == 738) begin
					state<=5;
					out<=198;
				end
				if(in == 739) begin
					state<=5;
					out<=199;
				end
				if(in == 740) begin
					state<=5;
					out<=200;
				end
				if(in == 741) begin
					state<=5;
					out<=201;
				end
				if(in == 742) begin
					state<=5;
					out<=202;
				end
				if(in == 743) begin
					state<=5;
					out<=203;
				end
				if(in == 744) begin
					state<=5;
					out<=204;
				end
				if(in == 745) begin
					state<=5;
					out<=205;
				end
				if(in == 746) begin
					state<=5;
					out<=206;
				end
				if(in == 747) begin
					state<=5;
					out<=207;
				end
				if(in == 748) begin
					state<=5;
					out<=208;
				end
				if(in == 749) begin
					state<=3;
					out<=209;
				end
				if(in == 750) begin
					state<=4;
					out<=210;
				end
				if(in == 751) begin
					state<=3;
					out<=211;
				end
				if(in == 752) begin
					state<=5;
					out<=212;
				end
				if(in == 753) begin
					state<=3;
					out<=213;
				end
				if(in == 754) begin
					state<=5;
					out<=214;
				end
				if(in == 755) begin
					state<=5;
					out<=215;
				end
				if(in == 756) begin
					state<=5;
					out<=216;
				end
				if(in == 757) begin
					state<=5;
					out<=217;
				end
				if(in == 758) begin
					state<=5;
					out<=218;
				end
				if(in == 759) begin
					state<=5;
					out<=219;
				end
				if(in == 760) begin
					state<=5;
					out<=220;
				end
				if(in == 761) begin
					state<=5;
					out<=221;
				end
				if(in == 762) begin
					state<=5;
					out<=222;
				end
				if(in == 763) begin
					state<=5;
					out<=223;
				end
				if(in == 764) begin
					state<=5;
					out<=224;
				end
				if(in == 765) begin
					state<=5;
					out<=225;
				end
				if(in == 766) begin
					state<=5;
					out<=226;
				end
				if(in == 767) begin
					state<=5;
					out<=227;
				end
				if(in == 768) begin
					state<=5;
					out<=228;
				end
				if(in == 769) begin
					state<=5;
					out<=229;
				end
				if(in == 770) begin
					state<=5;
					out<=230;
				end
				if(in == 771) begin
					state<=5;
					out<=231;
				end
				if(in == 772) begin
					state<=5;
					out<=232;
				end
				if(in == 773) begin
					state<=5;
					out<=233;
				end
				if(in == 774) begin
					state<=5;
					out<=234;
				end
				if(in == 775) begin
					state<=5;
					out<=235;
				end
				if(in == 776) begin
					state<=5;
					out<=236;
				end
				if(in == 777) begin
					state<=5;
					out<=237;
				end
				if(in == 778) begin
					state<=5;
					out<=238;
				end
				if(in == 779) begin
					state<=5;
					out<=239;
				end
				if(in == 780) begin
					state<=5;
					out<=240;
				end
				if(in == 781) begin
					state<=5;
					out<=241;
				end
				if(in == 782) begin
					state<=5;
					out<=242;
				end
				if(in == 783) begin
					state<=5;
					out<=243;
				end
				if(in == 784) begin
					state<=5;
					out<=244;
				end
				if(in == 785) begin
					state<=5;
					out<=245;
				end
				if(in == 786) begin
					state<=5;
					out<=246;
				end
				if(in == 787) begin
					state<=5;
					out<=247;
				end
				if(in == 788) begin
					state<=5;
					out<=248;
				end
				if(in == 789) begin
					state<=5;
					out<=249;
				end
				if(in == 790) begin
					state<=5;
					out<=250;
				end
				if(in == 791) begin
					state<=5;
					out<=251;
				end
				if(in == 792) begin
					state<=5;
					out<=252;
				end
				if(in == 793) begin
					state<=5;
					out<=253;
				end
				if(in == 794) begin
					state<=5;
					out<=254;
				end
				if(in == 795) begin
					state<=5;
					out<=255;
				end
				if(in == 796) begin
					state<=5;
					out<=0;
				end
				if(in == 797) begin
					state<=5;
					out<=1;
				end
				if(in == 798) begin
					state<=5;
					out<=2;
				end
				if(in == 799) begin
					state<=5;
					out<=3;
				end
				if(in == 800) begin
					state<=5;
					out<=4;
				end
				if(in == 801) begin
					state<=2;
					out<=5;
				end
				if(in == 802) begin
					state<=2;
					out<=6;
				end
				if(in == 803) begin
					state<=2;
					out<=7;
				end
				if(in == 804) begin
					state<=2;
					out<=8;
				end
				if(in == 805) begin
					state<=2;
					out<=9;
				end
				if(in == 806) begin
					state<=2;
					out<=10;
				end
				if(in == 807) begin
					state<=2;
					out<=11;
				end
				if(in == 808) begin
					state<=2;
					out<=12;
				end
				if(in == 809) begin
					state<=2;
					out<=13;
				end
				if(in == 810) begin
					state<=2;
					out<=14;
				end
				if(in == 811) begin
					state<=2;
					out<=15;
				end
				if(in == 812) begin
					state<=2;
					out<=16;
				end
				if(in == 813) begin
					state<=3;
					out<=17;
				end
				if(in == 814) begin
					state<=4;
					out<=18;
				end
				if(in == 815) begin
					state<=3;
					out<=19;
				end
				if(in == 816) begin
					state<=5;
					out<=20;
				end
				if(in == 817) begin
					state<=3;
					out<=21;
				end
				if(in == 818) begin
					state<=5;
					out<=22;
				end
				if(in == 819) begin
					state<=5;
					out<=23;
				end
				if(in == 820) begin
					state<=5;
					out<=24;
				end
				if(in == 821) begin
					state<=5;
					out<=25;
				end
				if(in == 822) begin
					state<=5;
					out<=26;
				end
				if(in == 823) begin
					state<=5;
					out<=27;
				end
				if(in == 824) begin
					state<=5;
					out<=28;
				end
				if(in == 825) begin
					state<=5;
					out<=29;
				end
				if(in == 826) begin
					state<=5;
					out<=30;
				end
				if(in == 827) begin
					state<=5;
					out<=31;
				end
				if(in == 828) begin
					state<=5;
					out<=32;
				end
				if(in == 829) begin
					state<=5;
					out<=33;
				end
				if(in == 830) begin
					state<=5;
					out<=34;
				end
				if(in == 831) begin
					state<=5;
					out<=35;
				end
				if(in == 832) begin
					state<=5;
					out<=36;
				end
				if(in == 833) begin
					state<=5;
					out<=37;
				end
				if(in == 834) begin
					state<=5;
					out<=38;
				end
				if(in == 835) begin
					state<=5;
					out<=39;
				end
				if(in == 836) begin
					state<=5;
					out<=40;
				end
				if(in == 837) begin
					state<=5;
					out<=41;
				end
				if(in == 838) begin
					state<=5;
					out<=42;
				end
				if(in == 839) begin
					state<=5;
					out<=43;
				end
				if(in == 840) begin
					state<=5;
					out<=44;
				end
				if(in == 841) begin
					state<=5;
					out<=45;
				end
				if(in == 842) begin
					state<=5;
					out<=46;
				end
				if(in == 843) begin
					state<=5;
					out<=47;
				end
				if(in == 844) begin
					state<=5;
					out<=48;
				end
				if(in == 845) begin
					state<=5;
					out<=49;
				end
				if(in == 846) begin
					state<=5;
					out<=50;
				end
				if(in == 847) begin
					state<=5;
					out<=51;
				end
				if(in == 848) begin
					state<=5;
					out<=52;
				end
				if(in == 849) begin
					state<=5;
					out<=53;
				end
				if(in == 850) begin
					state<=5;
					out<=54;
				end
				if(in == 851) begin
					state<=5;
					out<=55;
				end
				if(in == 852) begin
					state<=5;
					out<=56;
				end
				if(in == 853) begin
					state<=5;
					out<=57;
				end
				if(in == 854) begin
					state<=5;
					out<=58;
				end
				if(in == 855) begin
					state<=5;
					out<=59;
				end
				if(in == 856) begin
					state<=5;
					out<=60;
				end
				if(in == 857) begin
					state<=5;
					out<=61;
				end
				if(in == 858) begin
					state<=5;
					out<=62;
				end
				if(in == 859) begin
					state<=5;
					out<=63;
				end
				if(in == 860) begin
					state<=5;
					out<=64;
				end
				if(in == 861) begin
					state<=5;
					out<=65;
				end
				if(in == 862) begin
					state<=5;
					out<=66;
				end
				if(in == 863) begin
					state<=5;
					out<=67;
				end
				if(in == 864) begin
					state<=5;
					out<=68;
				end
				if(in == 865) begin
					state<=3;
					out<=69;
				end
				if(in == 866) begin
					state<=4;
					out<=70;
				end
				if(in == 867) begin
					state<=3;
					out<=71;
				end
				if(in == 868) begin
					state<=5;
					out<=72;
				end
				if(in == 869) begin
					state<=3;
					out<=73;
				end
				if(in == 870) begin
					state<=5;
					out<=74;
				end
				if(in == 871) begin
					state<=5;
					out<=75;
				end
				if(in == 872) begin
					state<=5;
					out<=76;
				end
				if(in == 873) begin
					state<=5;
					out<=77;
				end
				if(in == 874) begin
					state<=5;
					out<=78;
				end
				if(in == 875) begin
					state<=5;
					out<=79;
				end
				if(in == 876) begin
					state<=5;
					out<=80;
				end
				if(in == 877) begin
					state<=5;
					out<=81;
				end
				if(in == 878) begin
					state<=5;
					out<=82;
				end
				if(in == 879) begin
					state<=5;
					out<=83;
				end
				if(in == 880) begin
					state<=5;
					out<=84;
				end
				if(in == 881) begin
					state<=5;
					out<=85;
				end
				if(in == 882) begin
					state<=5;
					out<=86;
				end
				if(in == 883) begin
					state<=5;
					out<=87;
				end
				if(in == 884) begin
					state<=5;
					out<=88;
				end
				if(in == 885) begin
					state<=5;
					out<=89;
				end
				if(in == 886) begin
					state<=5;
					out<=90;
				end
				if(in == 887) begin
					state<=5;
					out<=91;
				end
				if(in == 888) begin
					state<=5;
					out<=92;
				end
				if(in == 889) begin
					state<=5;
					out<=93;
				end
				if(in == 890) begin
					state<=5;
					out<=94;
				end
				if(in == 891) begin
					state<=5;
					out<=95;
				end
				if(in == 892) begin
					state<=5;
					out<=96;
				end
				if(in == 893) begin
					state<=5;
					out<=97;
				end
				if(in == 894) begin
					state<=5;
					out<=98;
				end
				if(in == 895) begin
					state<=5;
					out<=99;
				end
				if(in == 896) begin
					state<=5;
					out<=100;
				end
				if(in == 897) begin
					state<=5;
					out<=101;
				end
				if(in == 898) begin
					state<=5;
					out<=102;
				end
				if(in == 899) begin
					state<=5;
					out<=103;
				end
				if(in == 900) begin
					state<=5;
					out<=104;
				end
				if(in == 901) begin
					state<=5;
					out<=105;
				end
				if(in == 902) begin
					state<=5;
					out<=106;
				end
				if(in == 903) begin
					state<=5;
					out<=107;
				end
				if(in == 904) begin
					state<=5;
					out<=108;
				end
				if(in == 905) begin
					state<=5;
					out<=109;
				end
				if(in == 906) begin
					state<=5;
					out<=110;
				end
				if(in == 907) begin
					state<=5;
					out<=111;
				end
				if(in == 908) begin
					state<=5;
					out<=112;
				end
				if(in == 909) begin
					state<=5;
					out<=113;
				end
				if(in == 910) begin
					state<=5;
					out<=114;
				end
				if(in == 911) begin
					state<=5;
					out<=115;
				end
				if(in == 912) begin
					state<=5;
					out<=116;
				end
				if(in == 913) begin
					state<=5;
					out<=117;
				end
				if(in == 914) begin
					state<=5;
					out<=118;
				end
				if(in == 915) begin
					state<=5;
					out<=119;
				end
				if(in == 916) begin
					state<=5;
					out<=120;
				end
				if(in == 917) begin
					state<=2;
					out<=121;
				end
				if(in == 918) begin
					state<=2;
					out<=122;
				end
				if(in == 919) begin
					state<=2;
					out<=123;
				end
				if(in == 920) begin
					state<=2;
					out<=124;
				end
				if(in == 921) begin
					state<=2;
					out<=125;
				end
				if(in == 922) begin
					state<=2;
					out<=126;
				end
				if(in == 923) begin
					state<=2;
					out<=127;
				end
				if(in == 924) begin
					state<=2;
					out<=128;
				end
				if(in == 925) begin
					state<=2;
					out<=129;
				end
				if(in == 926) begin
					state<=2;
					out<=130;
				end
				if(in == 927) begin
					state<=2;
					out<=131;
				end
				if(in == 928) begin
					state<=2;
					out<=132;
				end
			end
			5: begin
				if(in == 0) begin
					state<=3;
					out<=133;
				end
				if(in == 1) begin
					state<=1;
					out<=134;
				end
				if(in == 2) begin
					state<=5;
					out<=135;
				end
				if(in == 3) begin
					state<=3;
					out<=136;
				end
				if(in == 4) begin
					state<=5;
					out<=137;
				end
				if(in == 5) begin
					state<=3;
					out<=138;
				end
				if(in == 6) begin
					state<=5;
					out<=139;
				end
				if(in == 7) begin
					state<=5;
					out<=140;
				end
				if(in == 8) begin
					state<=5;
					out<=141;
				end
				if(in == 9) begin
					state<=5;
					out<=142;
				end
				if(in == 10) begin
					state<=5;
					out<=143;
				end
				if(in == 11) begin
					state<=5;
					out<=144;
				end
				if(in == 12) begin
					state<=5;
					out<=145;
				end
				if(in == 13) begin
					state<=5;
					out<=146;
				end
				if(in == 14) begin
					state<=5;
					out<=147;
				end
				if(in == 15) begin
					state<=5;
					out<=148;
				end
				if(in == 16) begin
					state<=5;
					out<=149;
				end
				if(in == 17) begin
					state<=5;
					out<=150;
				end
				if(in == 18) begin
					state<=5;
					out<=151;
				end
				if(in == 19) begin
					state<=5;
					out<=152;
				end
				if(in == 20) begin
					state<=5;
					out<=153;
				end
				if(in == 21) begin
					state<=6;
					out<=154;
				end
				if(in == 22) begin
					state<=6;
					out<=155;
				end
				if(in == 23) begin
					state<=6;
					out<=156;
				end
				if(in == 24) begin
					state<=6;
					out<=157;
				end
				if(in == 25) begin
					state<=6;
					out<=158;
				end
				if(in == 26) begin
					state<=6;
					out<=159;
				end
				if(in == 27) begin
					state<=6;
					out<=160;
				end
				if(in == 28) begin
					state<=6;
					out<=161;
				end
				if(in == 29) begin
					state<=6;
					out<=162;
				end
				if(in == 30) begin
					state<=6;
					out<=163;
				end
				if(in == 31) begin
					state<=6;
					out<=164;
				end
				if(in == 32) begin
					state<=6;
					out<=165;
				end
				if(in == 33) begin
					state<=6;
					out<=166;
				end
				if(in == 34) begin
					state<=6;
					out<=167;
				end
				if(in == 35) begin
					state<=6;
					out<=168;
				end
				if(in == 36) begin
					state<=6;
					out<=169;
				end
				if(in == 37) begin
					state<=5;
					out<=170;
				end
				if(in == 38) begin
					state<=5;
					out<=171;
				end
				if(in == 39) begin
					state<=5;
					out<=172;
				end
				if(in == 40) begin
					state<=5;
					out<=173;
				end
				if(in == 41) begin
					state<=5;
					out<=174;
				end
				if(in == 42) begin
					state<=5;
					out<=175;
				end
				if(in == 43) begin
					state<=5;
					out<=176;
				end
				if(in == 44) begin
					state<=5;
					out<=177;
				end
				if(in == 45) begin
					state<=5;
					out<=178;
				end
				if(in == 46) begin
					state<=5;
					out<=179;
				end
				if(in == 47) begin
					state<=5;
					out<=180;
				end
				if(in == 48) begin
					state<=5;
					out<=181;
				end
				if(in == 49) begin
					state<=5;
					out<=182;
				end
				if(in == 50) begin
					state<=5;
					out<=183;
				end
				if(in == 51) begin
					state<=5;
					out<=184;
				end
				if(in == 52) begin
					state<=5;
					out<=185;
				end
				if(in == 53) begin
					state<=3;
					out<=186;
				end
				if(in == 54) begin
					state<=5;
					out<=187;
				end
				if(in == 55) begin
					state<=3;
					out<=188;
				end
				if(in == 56) begin
					state<=5;
					out<=189;
				end
				if(in == 57) begin
					state<=3;
					out<=190;
				end
				if(in == 58) begin
					state<=5;
					out<=191;
				end
				if(in == 59) begin
					state<=5;
					out<=192;
				end
				if(in == 60) begin
					state<=5;
					out<=193;
				end
				if(in == 61) begin
					state<=5;
					out<=194;
				end
				if(in == 62) begin
					state<=5;
					out<=195;
				end
				if(in == 63) begin
					state<=5;
					out<=196;
				end
				if(in == 64) begin
					state<=5;
					out<=197;
				end
				if(in == 65) begin
					state<=5;
					out<=198;
				end
				if(in == 66) begin
					state<=5;
					out<=199;
				end
				if(in == 67) begin
					state<=5;
					out<=200;
				end
				if(in == 68) begin
					state<=5;
					out<=201;
				end
				if(in == 69) begin
					state<=5;
					out<=202;
				end
				if(in == 70) begin
					state<=5;
					out<=203;
				end
				if(in == 71) begin
					state<=5;
					out<=204;
				end
				if(in == 72) begin
					state<=5;
					out<=205;
				end
				if(in == 73) begin
					state<=6;
					out<=206;
				end
				if(in == 74) begin
					state<=6;
					out<=207;
				end
				if(in == 75) begin
					state<=6;
					out<=208;
				end
				if(in == 76) begin
					state<=6;
					out<=209;
				end
				if(in == 77) begin
					state<=6;
					out<=210;
				end
				if(in == 78) begin
					state<=6;
					out<=211;
				end
				if(in == 79) begin
					state<=6;
					out<=212;
				end
				if(in == 80) begin
					state<=6;
					out<=213;
				end
				if(in == 81) begin
					state<=6;
					out<=214;
				end
				if(in == 82) begin
					state<=6;
					out<=215;
				end
				if(in == 83) begin
					state<=6;
					out<=216;
				end
				if(in == 84) begin
					state<=6;
					out<=217;
				end
				if(in == 85) begin
					state<=6;
					out<=218;
				end
				if(in == 86) begin
					state<=6;
					out<=219;
				end
				if(in == 87) begin
					state<=6;
					out<=220;
				end
				if(in == 88) begin
					state<=6;
					out<=221;
				end
				if(in == 89) begin
					state<=5;
					out<=222;
				end
				if(in == 90) begin
					state<=5;
					out<=223;
				end
				if(in == 91) begin
					state<=5;
					out<=224;
				end
				if(in == 92) begin
					state<=5;
					out<=225;
				end
				if(in == 93) begin
					state<=5;
					out<=226;
				end
				if(in == 94) begin
					state<=5;
					out<=227;
				end
				if(in == 95) begin
					state<=5;
					out<=228;
				end
				if(in == 96) begin
					state<=5;
					out<=229;
				end
				if(in == 97) begin
					state<=5;
					out<=230;
				end
				if(in == 98) begin
					state<=5;
					out<=231;
				end
				if(in == 99) begin
					state<=5;
					out<=232;
				end
				if(in == 100) begin
					state<=5;
					out<=233;
				end
				if(in == 101) begin
					state<=5;
					out<=234;
				end
				if(in == 102) begin
					state<=5;
					out<=235;
				end
				if(in == 103) begin
					state<=5;
					out<=236;
				end
				if(in == 104) begin
					state<=5;
					out<=237;
				end
				if(in == 105) begin
					state<=2;
					out<=238;
				end
				if(in == 106) begin
					state<=2;
					out<=239;
				end
				if(in == 107) begin
					state<=2;
					out<=240;
				end
				if(in == 108) begin
					state<=2;
					out<=241;
				end
				if(in == 109) begin
					state<=2;
					out<=242;
				end
				if(in == 110) begin
					state<=2;
					out<=243;
				end
				if(in == 111) begin
					state<=2;
					out<=244;
				end
				if(in == 112) begin
					state<=2;
					out<=245;
				end
				if(in == 113) begin
					state<=2;
					out<=246;
				end
				if(in == 114) begin
					state<=2;
					out<=247;
				end
				if(in == 115) begin
					state<=2;
					out<=248;
				end
				if(in == 116) begin
					state<=2;
					out<=249;
				end
				if(in == 117) begin
					state<=3;
					out<=250;
				end
				if(in == 118) begin
					state<=5;
					out<=251;
				end
				if(in == 119) begin
					state<=3;
					out<=252;
				end
				if(in == 120) begin
					state<=5;
					out<=253;
				end
				if(in == 121) begin
					state<=3;
					out<=254;
				end
				if(in == 122) begin
					state<=5;
					out<=255;
				end
				if(in == 123) begin
					state<=5;
					out<=0;
				end
				if(in == 124) begin
					state<=5;
					out<=1;
				end
				if(in == 125) begin
					state<=5;
					out<=2;
				end
				if(in == 126) begin
					state<=5;
					out<=3;
				end
				if(in == 127) begin
					state<=5;
					out<=4;
				end
				if(in == 128) begin
					state<=5;
					out<=5;
				end
				if(in == 129) begin
					state<=5;
					out<=6;
				end
				if(in == 130) begin
					state<=5;
					out<=7;
				end
				if(in == 131) begin
					state<=5;
					out<=8;
				end
				if(in == 132) begin
					state<=5;
					out<=9;
				end
				if(in == 133) begin
					state<=5;
					out<=10;
				end
				if(in == 134) begin
					state<=5;
					out<=11;
				end
				if(in == 135) begin
					state<=5;
					out<=12;
				end
				if(in == 136) begin
					state<=5;
					out<=13;
				end
				if(in == 137) begin
					state<=6;
					out<=14;
				end
				if(in == 138) begin
					state<=6;
					out<=15;
				end
				if(in == 139) begin
					state<=6;
					out<=16;
				end
				if(in == 140) begin
					state<=6;
					out<=17;
				end
				if(in == 141) begin
					state<=6;
					out<=18;
				end
				if(in == 142) begin
					state<=6;
					out<=19;
				end
				if(in == 143) begin
					state<=6;
					out<=20;
				end
				if(in == 144) begin
					state<=6;
					out<=21;
				end
				if(in == 145) begin
					state<=6;
					out<=22;
				end
				if(in == 146) begin
					state<=6;
					out<=23;
				end
				if(in == 147) begin
					state<=6;
					out<=24;
				end
				if(in == 148) begin
					state<=6;
					out<=25;
				end
				if(in == 149) begin
					state<=6;
					out<=26;
				end
				if(in == 150) begin
					state<=6;
					out<=27;
				end
				if(in == 151) begin
					state<=6;
					out<=28;
				end
				if(in == 152) begin
					state<=6;
					out<=29;
				end
				if(in == 153) begin
					state<=5;
					out<=30;
				end
				if(in == 154) begin
					state<=5;
					out<=31;
				end
				if(in == 155) begin
					state<=5;
					out<=32;
				end
				if(in == 156) begin
					state<=5;
					out<=33;
				end
				if(in == 157) begin
					state<=5;
					out<=34;
				end
				if(in == 158) begin
					state<=5;
					out<=35;
				end
				if(in == 159) begin
					state<=5;
					out<=36;
				end
				if(in == 160) begin
					state<=5;
					out<=37;
				end
				if(in == 161) begin
					state<=5;
					out<=38;
				end
				if(in == 162) begin
					state<=5;
					out<=39;
				end
				if(in == 163) begin
					state<=5;
					out<=40;
				end
				if(in == 164) begin
					state<=5;
					out<=41;
				end
				if(in == 165) begin
					state<=5;
					out<=42;
				end
				if(in == 166) begin
					state<=5;
					out<=43;
				end
				if(in == 167) begin
					state<=5;
					out<=44;
				end
				if(in == 168) begin
					state<=5;
					out<=45;
				end
				if(in == 169) begin
					state<=3;
					out<=46;
				end
				if(in == 170) begin
					state<=5;
					out<=47;
				end
				if(in == 171) begin
					state<=3;
					out<=48;
				end
				if(in == 172) begin
					state<=5;
					out<=49;
				end
				if(in == 173) begin
					state<=3;
					out<=50;
				end
				if(in == 174) begin
					state<=5;
					out<=51;
				end
				if(in == 175) begin
					state<=5;
					out<=52;
				end
				if(in == 176) begin
					state<=5;
					out<=53;
				end
				if(in == 177) begin
					state<=5;
					out<=54;
				end
				if(in == 178) begin
					state<=5;
					out<=55;
				end
				if(in == 179) begin
					state<=5;
					out<=56;
				end
				if(in == 180) begin
					state<=5;
					out<=57;
				end
				if(in == 181) begin
					state<=5;
					out<=58;
				end
				if(in == 182) begin
					state<=5;
					out<=59;
				end
				if(in == 183) begin
					state<=5;
					out<=60;
				end
				if(in == 184) begin
					state<=5;
					out<=61;
				end
				if(in == 185) begin
					state<=5;
					out<=62;
				end
				if(in == 186) begin
					state<=5;
					out<=63;
				end
				if(in == 187) begin
					state<=5;
					out<=64;
				end
				if(in == 188) begin
					state<=5;
					out<=65;
				end
				if(in == 189) begin
					state<=6;
					out<=66;
				end
				if(in == 190) begin
					state<=6;
					out<=67;
				end
				if(in == 191) begin
					state<=6;
					out<=68;
				end
				if(in == 192) begin
					state<=6;
					out<=69;
				end
				if(in == 193) begin
					state<=6;
					out<=70;
				end
				if(in == 194) begin
					state<=6;
					out<=71;
				end
				if(in == 195) begin
					state<=6;
					out<=72;
				end
				if(in == 196) begin
					state<=6;
					out<=73;
				end
				if(in == 197) begin
					state<=6;
					out<=74;
				end
				if(in == 198) begin
					state<=6;
					out<=75;
				end
				if(in == 199) begin
					state<=6;
					out<=76;
				end
				if(in == 200) begin
					state<=6;
					out<=77;
				end
				if(in == 201) begin
					state<=6;
					out<=78;
				end
				if(in == 202) begin
					state<=6;
					out<=79;
				end
				if(in == 203) begin
					state<=6;
					out<=80;
				end
				if(in == 204) begin
					state<=6;
					out<=81;
				end
				if(in == 205) begin
					state<=5;
					out<=82;
				end
				if(in == 206) begin
					state<=5;
					out<=83;
				end
				if(in == 207) begin
					state<=5;
					out<=84;
				end
				if(in == 208) begin
					state<=5;
					out<=85;
				end
				if(in == 209) begin
					state<=5;
					out<=86;
				end
				if(in == 210) begin
					state<=5;
					out<=87;
				end
				if(in == 211) begin
					state<=5;
					out<=88;
				end
				if(in == 212) begin
					state<=5;
					out<=89;
				end
				if(in == 213) begin
					state<=5;
					out<=90;
				end
				if(in == 214) begin
					state<=5;
					out<=91;
				end
				if(in == 215) begin
					state<=5;
					out<=92;
				end
				if(in == 216) begin
					state<=5;
					out<=93;
				end
				if(in == 217) begin
					state<=5;
					out<=94;
				end
				if(in == 218) begin
					state<=5;
					out<=95;
				end
				if(in == 219) begin
					state<=5;
					out<=96;
				end
				if(in == 220) begin
					state<=5;
					out<=97;
				end
				if(in == 221) begin
					state<=2;
					out<=98;
				end
				if(in == 222) begin
					state<=2;
					out<=99;
				end
				if(in == 223) begin
					state<=2;
					out<=100;
				end
				if(in == 224) begin
					state<=2;
					out<=101;
				end
				if(in == 225) begin
					state<=2;
					out<=102;
				end
				if(in == 226) begin
					state<=2;
					out<=103;
				end
				if(in == 227) begin
					state<=2;
					out<=104;
				end
				if(in == 228) begin
					state<=2;
					out<=105;
				end
				if(in == 229) begin
					state<=2;
					out<=106;
				end
				if(in == 230) begin
					state<=2;
					out<=107;
				end
				if(in == 231) begin
					state<=2;
					out<=108;
				end
				if(in == 232) begin
					state<=2;
					out<=109;
				end
				if(in == 233) begin
					state<=3;
					out<=110;
				end
				if(in == 234) begin
					state<=5;
					out<=111;
				end
				if(in == 235) begin
					state<=3;
					out<=112;
				end
				if(in == 236) begin
					state<=5;
					out<=113;
				end
				if(in == 237) begin
					state<=3;
					out<=114;
				end
				if(in == 238) begin
					state<=5;
					out<=115;
				end
				if(in == 239) begin
					state<=5;
					out<=116;
				end
				if(in == 240) begin
					state<=5;
					out<=117;
				end
				if(in == 241) begin
					state<=5;
					out<=118;
				end
				if(in == 242) begin
					state<=5;
					out<=119;
				end
				if(in == 243) begin
					state<=5;
					out<=120;
				end
				if(in == 244) begin
					state<=5;
					out<=121;
				end
				if(in == 245) begin
					state<=5;
					out<=122;
				end
				if(in == 246) begin
					state<=5;
					out<=123;
				end
				if(in == 247) begin
					state<=5;
					out<=124;
				end
				if(in == 248) begin
					state<=5;
					out<=125;
				end
				if(in == 249) begin
					state<=5;
					out<=126;
				end
				if(in == 250) begin
					state<=5;
					out<=127;
				end
				if(in == 251) begin
					state<=5;
					out<=128;
				end
				if(in == 252) begin
					state<=5;
					out<=129;
				end
				if(in == 253) begin
					state<=6;
					out<=130;
				end
				if(in == 254) begin
					state<=6;
					out<=131;
				end
				if(in == 255) begin
					state<=6;
					out<=132;
				end
				if(in == 256) begin
					state<=6;
					out<=133;
				end
				if(in == 257) begin
					state<=6;
					out<=134;
				end
				if(in == 258) begin
					state<=6;
					out<=135;
				end
				if(in == 259) begin
					state<=6;
					out<=136;
				end
				if(in == 260) begin
					state<=6;
					out<=137;
				end
				if(in == 261) begin
					state<=6;
					out<=138;
				end
				if(in == 262) begin
					state<=6;
					out<=139;
				end
				if(in == 263) begin
					state<=6;
					out<=140;
				end
				if(in == 264) begin
					state<=6;
					out<=141;
				end
				if(in == 265) begin
					state<=6;
					out<=142;
				end
				if(in == 266) begin
					state<=6;
					out<=143;
				end
				if(in == 267) begin
					state<=6;
					out<=144;
				end
				if(in == 268) begin
					state<=6;
					out<=145;
				end
				if(in == 269) begin
					state<=5;
					out<=146;
				end
				if(in == 270) begin
					state<=5;
					out<=147;
				end
				if(in == 271) begin
					state<=5;
					out<=148;
				end
				if(in == 272) begin
					state<=5;
					out<=149;
				end
				if(in == 273) begin
					state<=5;
					out<=150;
				end
				if(in == 274) begin
					state<=5;
					out<=151;
				end
				if(in == 275) begin
					state<=5;
					out<=152;
				end
				if(in == 276) begin
					state<=5;
					out<=153;
				end
				if(in == 277) begin
					state<=5;
					out<=154;
				end
				if(in == 278) begin
					state<=5;
					out<=155;
				end
				if(in == 279) begin
					state<=5;
					out<=156;
				end
				if(in == 280) begin
					state<=5;
					out<=157;
				end
				if(in == 281) begin
					state<=5;
					out<=158;
				end
				if(in == 282) begin
					state<=5;
					out<=159;
				end
				if(in == 283) begin
					state<=5;
					out<=160;
				end
				if(in == 284) begin
					state<=5;
					out<=161;
				end
				if(in == 285) begin
					state<=3;
					out<=162;
				end
				if(in == 286) begin
					state<=5;
					out<=163;
				end
				if(in == 287) begin
					state<=3;
					out<=164;
				end
				if(in == 288) begin
					state<=5;
					out<=165;
				end
				if(in == 289) begin
					state<=3;
					out<=166;
				end
				if(in == 290) begin
					state<=5;
					out<=167;
				end
				if(in == 291) begin
					state<=5;
					out<=168;
				end
				if(in == 292) begin
					state<=5;
					out<=169;
				end
				if(in == 293) begin
					state<=5;
					out<=170;
				end
				if(in == 294) begin
					state<=5;
					out<=171;
				end
				if(in == 295) begin
					state<=5;
					out<=172;
				end
				if(in == 296) begin
					state<=5;
					out<=173;
				end
				if(in == 297) begin
					state<=5;
					out<=174;
				end
				if(in == 298) begin
					state<=5;
					out<=175;
				end
				if(in == 299) begin
					state<=5;
					out<=176;
				end
				if(in == 300) begin
					state<=5;
					out<=177;
				end
				if(in == 301) begin
					state<=5;
					out<=178;
				end
				if(in == 302) begin
					state<=5;
					out<=179;
				end
				if(in == 303) begin
					state<=5;
					out<=180;
				end
				if(in == 304) begin
					state<=5;
					out<=181;
				end
				if(in == 305) begin
					state<=6;
					out<=182;
				end
				if(in == 306) begin
					state<=6;
					out<=183;
				end
				if(in == 307) begin
					state<=6;
					out<=184;
				end
				if(in == 308) begin
					state<=6;
					out<=185;
				end
				if(in == 309) begin
					state<=6;
					out<=186;
				end
				if(in == 310) begin
					state<=6;
					out<=187;
				end
				if(in == 311) begin
					state<=6;
					out<=188;
				end
				if(in == 312) begin
					state<=6;
					out<=189;
				end
				if(in == 313) begin
					state<=6;
					out<=190;
				end
				if(in == 314) begin
					state<=6;
					out<=191;
				end
				if(in == 315) begin
					state<=6;
					out<=192;
				end
				if(in == 316) begin
					state<=6;
					out<=193;
				end
				if(in == 317) begin
					state<=6;
					out<=194;
				end
				if(in == 318) begin
					state<=6;
					out<=195;
				end
				if(in == 319) begin
					state<=6;
					out<=196;
				end
				if(in == 320) begin
					state<=6;
					out<=197;
				end
				if(in == 321) begin
					state<=5;
					out<=198;
				end
				if(in == 322) begin
					state<=5;
					out<=199;
				end
				if(in == 323) begin
					state<=5;
					out<=200;
				end
				if(in == 324) begin
					state<=5;
					out<=201;
				end
				if(in == 325) begin
					state<=5;
					out<=202;
				end
				if(in == 326) begin
					state<=5;
					out<=203;
				end
				if(in == 327) begin
					state<=5;
					out<=204;
				end
				if(in == 328) begin
					state<=5;
					out<=205;
				end
				if(in == 329) begin
					state<=5;
					out<=206;
				end
				if(in == 330) begin
					state<=5;
					out<=207;
				end
				if(in == 331) begin
					state<=5;
					out<=208;
				end
				if(in == 332) begin
					state<=5;
					out<=209;
				end
				if(in == 333) begin
					state<=5;
					out<=210;
				end
				if(in == 334) begin
					state<=5;
					out<=211;
				end
				if(in == 335) begin
					state<=5;
					out<=212;
				end
				if(in == 336) begin
					state<=5;
					out<=213;
				end
				if(in == 337) begin
					state<=2;
					out<=214;
				end
				if(in == 338) begin
					state<=2;
					out<=215;
				end
				if(in == 339) begin
					state<=2;
					out<=216;
				end
				if(in == 340) begin
					state<=2;
					out<=217;
				end
				if(in == 341) begin
					state<=2;
					out<=218;
				end
				if(in == 342) begin
					state<=2;
					out<=219;
				end
				if(in == 343) begin
					state<=2;
					out<=220;
				end
				if(in == 344) begin
					state<=2;
					out<=221;
				end
				if(in == 345) begin
					state<=2;
					out<=222;
				end
				if(in == 346) begin
					state<=2;
					out<=223;
				end
				if(in == 347) begin
					state<=2;
					out<=224;
				end
				if(in == 348) begin
					state<=2;
					out<=225;
				end
				if(in == 349) begin
					state<=3;
					out<=226;
				end
				if(in == 350) begin
					state<=5;
					out<=227;
				end
				if(in == 351) begin
					state<=3;
					out<=228;
				end
				if(in == 352) begin
					state<=5;
					out<=229;
				end
				if(in == 353) begin
					state<=3;
					out<=230;
				end
				if(in == 354) begin
					state<=5;
					out<=231;
				end
				if(in == 355) begin
					state<=5;
					out<=232;
				end
				if(in == 356) begin
					state<=5;
					out<=233;
				end
				if(in == 357) begin
					state<=5;
					out<=234;
				end
				if(in == 358) begin
					state<=5;
					out<=235;
				end
				if(in == 359) begin
					state<=5;
					out<=236;
				end
				if(in == 360) begin
					state<=5;
					out<=237;
				end
				if(in == 361) begin
					state<=5;
					out<=238;
				end
				if(in == 362) begin
					state<=5;
					out<=239;
				end
				if(in == 363) begin
					state<=5;
					out<=240;
				end
				if(in == 364) begin
					state<=5;
					out<=241;
				end
				if(in == 365) begin
					state<=5;
					out<=242;
				end
				if(in == 366) begin
					state<=5;
					out<=243;
				end
				if(in == 367) begin
					state<=5;
					out<=244;
				end
				if(in == 368) begin
					state<=5;
					out<=245;
				end
				if(in == 369) begin
					state<=6;
					out<=246;
				end
				if(in == 370) begin
					state<=6;
					out<=247;
				end
				if(in == 371) begin
					state<=6;
					out<=248;
				end
				if(in == 372) begin
					state<=6;
					out<=249;
				end
				if(in == 373) begin
					state<=6;
					out<=250;
				end
				if(in == 374) begin
					state<=6;
					out<=251;
				end
				if(in == 375) begin
					state<=6;
					out<=252;
				end
				if(in == 376) begin
					state<=6;
					out<=253;
				end
				if(in == 377) begin
					state<=6;
					out<=254;
				end
				if(in == 378) begin
					state<=6;
					out<=255;
				end
				if(in == 379) begin
					state<=6;
					out<=0;
				end
				if(in == 380) begin
					state<=6;
					out<=1;
				end
				if(in == 381) begin
					state<=6;
					out<=2;
				end
				if(in == 382) begin
					state<=6;
					out<=3;
				end
				if(in == 383) begin
					state<=6;
					out<=4;
				end
				if(in == 384) begin
					state<=6;
					out<=5;
				end
				if(in == 385) begin
					state<=5;
					out<=6;
				end
				if(in == 386) begin
					state<=5;
					out<=7;
				end
				if(in == 387) begin
					state<=5;
					out<=8;
				end
				if(in == 388) begin
					state<=5;
					out<=9;
				end
				if(in == 389) begin
					state<=5;
					out<=10;
				end
				if(in == 390) begin
					state<=5;
					out<=11;
				end
				if(in == 391) begin
					state<=5;
					out<=12;
				end
				if(in == 392) begin
					state<=5;
					out<=13;
				end
				if(in == 393) begin
					state<=5;
					out<=14;
				end
				if(in == 394) begin
					state<=5;
					out<=15;
				end
				if(in == 395) begin
					state<=5;
					out<=16;
				end
				if(in == 396) begin
					state<=5;
					out<=17;
				end
				if(in == 397) begin
					state<=5;
					out<=18;
				end
				if(in == 398) begin
					state<=5;
					out<=19;
				end
				if(in == 399) begin
					state<=5;
					out<=20;
				end
				if(in == 400) begin
					state<=5;
					out<=21;
				end
				if(in == 401) begin
					state<=3;
					out<=22;
				end
				if(in == 402) begin
					state<=5;
					out<=23;
				end
				if(in == 403) begin
					state<=3;
					out<=24;
				end
				if(in == 404) begin
					state<=5;
					out<=25;
				end
				if(in == 405) begin
					state<=3;
					out<=26;
				end
				if(in == 406) begin
					state<=5;
					out<=27;
				end
				if(in == 407) begin
					state<=5;
					out<=28;
				end
				if(in == 408) begin
					state<=5;
					out<=29;
				end
				if(in == 409) begin
					state<=5;
					out<=30;
				end
				if(in == 410) begin
					state<=5;
					out<=31;
				end
				if(in == 411) begin
					state<=5;
					out<=32;
				end
				if(in == 412) begin
					state<=5;
					out<=33;
				end
				if(in == 413) begin
					state<=5;
					out<=34;
				end
				if(in == 414) begin
					state<=5;
					out<=35;
				end
				if(in == 415) begin
					state<=5;
					out<=36;
				end
				if(in == 416) begin
					state<=5;
					out<=37;
				end
				if(in == 417) begin
					state<=5;
					out<=38;
				end
				if(in == 418) begin
					state<=5;
					out<=39;
				end
				if(in == 419) begin
					state<=5;
					out<=40;
				end
				if(in == 420) begin
					state<=5;
					out<=41;
				end
				if(in == 421) begin
					state<=6;
					out<=42;
				end
				if(in == 422) begin
					state<=6;
					out<=43;
				end
				if(in == 423) begin
					state<=6;
					out<=44;
				end
				if(in == 424) begin
					state<=6;
					out<=45;
				end
				if(in == 425) begin
					state<=6;
					out<=46;
				end
				if(in == 426) begin
					state<=6;
					out<=47;
				end
				if(in == 427) begin
					state<=6;
					out<=48;
				end
				if(in == 428) begin
					state<=6;
					out<=49;
				end
				if(in == 429) begin
					state<=6;
					out<=50;
				end
				if(in == 430) begin
					state<=6;
					out<=51;
				end
				if(in == 431) begin
					state<=6;
					out<=52;
				end
				if(in == 432) begin
					state<=6;
					out<=53;
				end
				if(in == 433) begin
					state<=6;
					out<=54;
				end
				if(in == 434) begin
					state<=6;
					out<=55;
				end
				if(in == 435) begin
					state<=6;
					out<=56;
				end
				if(in == 436) begin
					state<=6;
					out<=57;
				end
				if(in == 437) begin
					state<=5;
					out<=58;
				end
				if(in == 438) begin
					state<=5;
					out<=59;
				end
				if(in == 439) begin
					state<=5;
					out<=60;
				end
				if(in == 440) begin
					state<=5;
					out<=61;
				end
				if(in == 441) begin
					state<=5;
					out<=62;
				end
				if(in == 442) begin
					state<=5;
					out<=63;
				end
				if(in == 443) begin
					state<=5;
					out<=64;
				end
				if(in == 444) begin
					state<=5;
					out<=65;
				end
				if(in == 445) begin
					state<=5;
					out<=66;
				end
				if(in == 446) begin
					state<=5;
					out<=67;
				end
				if(in == 447) begin
					state<=5;
					out<=68;
				end
				if(in == 448) begin
					state<=5;
					out<=69;
				end
				if(in == 449) begin
					state<=5;
					out<=70;
				end
				if(in == 450) begin
					state<=5;
					out<=71;
				end
				if(in == 451) begin
					state<=5;
					out<=72;
				end
				if(in == 452) begin
					state<=5;
					out<=73;
				end
				if(in == 453) begin
					state<=2;
					out<=74;
				end
				if(in == 454) begin
					state<=2;
					out<=75;
				end
				if(in == 455) begin
					state<=2;
					out<=76;
				end
				if(in == 456) begin
					state<=2;
					out<=77;
				end
				if(in == 457) begin
					state<=2;
					out<=78;
				end
				if(in == 458) begin
					state<=2;
					out<=79;
				end
				if(in == 459) begin
					state<=2;
					out<=80;
				end
				if(in == 460) begin
					state<=2;
					out<=81;
				end
				if(in == 461) begin
					state<=2;
					out<=82;
				end
				if(in == 462) begin
					state<=2;
					out<=83;
				end
				if(in == 463) begin
					state<=2;
					out<=84;
				end
				if(in == 464) begin
					state<=2;
					out<=85;
				end
				if(in == 465) begin
					state<=3;
					out<=86;
				end
				if(in == 466) begin
					state<=5;
					out<=87;
				end
				if(in == 467) begin
					state<=3;
					out<=88;
				end
				if(in == 468) begin
					state<=5;
					out<=89;
				end
				if(in == 469) begin
					state<=3;
					out<=90;
				end
				if(in == 470) begin
					state<=5;
					out<=91;
				end
				if(in == 471) begin
					state<=5;
					out<=92;
				end
				if(in == 472) begin
					state<=5;
					out<=93;
				end
				if(in == 473) begin
					state<=5;
					out<=94;
				end
				if(in == 474) begin
					state<=5;
					out<=95;
				end
				if(in == 475) begin
					state<=5;
					out<=96;
				end
				if(in == 476) begin
					state<=5;
					out<=97;
				end
				if(in == 477) begin
					state<=5;
					out<=98;
				end
				if(in == 478) begin
					state<=5;
					out<=99;
				end
				if(in == 479) begin
					state<=5;
					out<=100;
				end
				if(in == 480) begin
					state<=5;
					out<=101;
				end
				if(in == 481) begin
					state<=5;
					out<=102;
				end
				if(in == 482) begin
					state<=5;
					out<=103;
				end
				if(in == 483) begin
					state<=5;
					out<=104;
				end
				if(in == 484) begin
					state<=5;
					out<=105;
				end
				if(in == 485) begin
					state<=6;
					out<=106;
				end
				if(in == 486) begin
					state<=6;
					out<=107;
				end
				if(in == 487) begin
					state<=6;
					out<=108;
				end
				if(in == 488) begin
					state<=6;
					out<=109;
				end
				if(in == 489) begin
					state<=6;
					out<=110;
				end
				if(in == 490) begin
					state<=6;
					out<=111;
				end
				if(in == 491) begin
					state<=6;
					out<=112;
				end
				if(in == 492) begin
					state<=6;
					out<=113;
				end
				if(in == 493) begin
					state<=6;
					out<=114;
				end
				if(in == 494) begin
					state<=6;
					out<=115;
				end
				if(in == 495) begin
					state<=6;
					out<=116;
				end
				if(in == 496) begin
					state<=6;
					out<=117;
				end
				if(in == 497) begin
					state<=6;
					out<=118;
				end
				if(in == 498) begin
					state<=6;
					out<=119;
				end
				if(in == 499) begin
					state<=6;
					out<=120;
				end
				if(in == 500) begin
					state<=6;
					out<=121;
				end
				if(in == 501) begin
					state<=5;
					out<=122;
				end
				if(in == 502) begin
					state<=5;
					out<=123;
				end
				if(in == 503) begin
					state<=5;
					out<=124;
				end
				if(in == 504) begin
					state<=5;
					out<=125;
				end
				if(in == 505) begin
					state<=5;
					out<=126;
				end
				if(in == 506) begin
					state<=5;
					out<=127;
				end
				if(in == 507) begin
					state<=5;
					out<=128;
				end
				if(in == 508) begin
					state<=5;
					out<=129;
				end
				if(in == 509) begin
					state<=5;
					out<=130;
				end
				if(in == 510) begin
					state<=5;
					out<=131;
				end
				if(in == 511) begin
					state<=5;
					out<=132;
				end
				if(in == 512) begin
					state<=5;
					out<=133;
				end
				if(in == 513) begin
					state<=5;
					out<=134;
				end
				if(in == 514) begin
					state<=5;
					out<=135;
				end
				if(in == 515) begin
					state<=5;
					out<=136;
				end
				if(in == 516) begin
					state<=5;
					out<=137;
				end
				if(in == 517) begin
					state<=3;
					out<=138;
				end
				if(in == 518) begin
					state<=5;
					out<=139;
				end
				if(in == 519) begin
					state<=3;
					out<=140;
				end
				if(in == 520) begin
					state<=5;
					out<=141;
				end
				if(in == 521) begin
					state<=3;
					out<=142;
				end
				if(in == 522) begin
					state<=5;
					out<=143;
				end
				if(in == 523) begin
					state<=5;
					out<=144;
				end
				if(in == 524) begin
					state<=5;
					out<=145;
				end
				if(in == 525) begin
					state<=5;
					out<=146;
				end
				if(in == 526) begin
					state<=5;
					out<=147;
				end
				if(in == 527) begin
					state<=5;
					out<=148;
				end
				if(in == 528) begin
					state<=5;
					out<=149;
				end
				if(in == 529) begin
					state<=5;
					out<=150;
				end
				if(in == 530) begin
					state<=5;
					out<=151;
				end
				if(in == 531) begin
					state<=5;
					out<=152;
				end
				if(in == 532) begin
					state<=5;
					out<=153;
				end
				if(in == 533) begin
					state<=5;
					out<=154;
				end
				if(in == 534) begin
					state<=5;
					out<=155;
				end
				if(in == 535) begin
					state<=5;
					out<=156;
				end
				if(in == 536) begin
					state<=5;
					out<=157;
				end
				if(in == 537) begin
					state<=6;
					out<=158;
				end
				if(in == 538) begin
					state<=6;
					out<=159;
				end
				if(in == 539) begin
					state<=6;
					out<=160;
				end
				if(in == 540) begin
					state<=6;
					out<=161;
				end
				if(in == 541) begin
					state<=6;
					out<=162;
				end
				if(in == 542) begin
					state<=6;
					out<=163;
				end
				if(in == 543) begin
					state<=6;
					out<=164;
				end
				if(in == 544) begin
					state<=6;
					out<=165;
				end
				if(in == 545) begin
					state<=6;
					out<=166;
				end
				if(in == 546) begin
					state<=6;
					out<=167;
				end
				if(in == 547) begin
					state<=6;
					out<=168;
				end
				if(in == 548) begin
					state<=6;
					out<=169;
				end
				if(in == 549) begin
					state<=6;
					out<=170;
				end
				if(in == 550) begin
					state<=6;
					out<=171;
				end
				if(in == 551) begin
					state<=6;
					out<=172;
				end
				if(in == 552) begin
					state<=6;
					out<=173;
				end
				if(in == 553) begin
					state<=5;
					out<=174;
				end
				if(in == 554) begin
					state<=5;
					out<=175;
				end
				if(in == 555) begin
					state<=5;
					out<=176;
				end
				if(in == 556) begin
					state<=5;
					out<=177;
				end
				if(in == 557) begin
					state<=5;
					out<=178;
				end
				if(in == 558) begin
					state<=5;
					out<=179;
				end
				if(in == 559) begin
					state<=5;
					out<=180;
				end
				if(in == 560) begin
					state<=5;
					out<=181;
				end
				if(in == 561) begin
					state<=5;
					out<=182;
				end
				if(in == 562) begin
					state<=5;
					out<=183;
				end
				if(in == 563) begin
					state<=5;
					out<=184;
				end
				if(in == 564) begin
					state<=5;
					out<=185;
				end
				if(in == 565) begin
					state<=5;
					out<=186;
				end
				if(in == 566) begin
					state<=5;
					out<=187;
				end
				if(in == 567) begin
					state<=5;
					out<=188;
				end
				if(in == 568) begin
					state<=5;
					out<=189;
				end
				if(in == 569) begin
					state<=2;
					out<=190;
				end
				if(in == 570) begin
					state<=2;
					out<=191;
				end
				if(in == 571) begin
					state<=2;
					out<=192;
				end
				if(in == 572) begin
					state<=2;
					out<=193;
				end
				if(in == 573) begin
					state<=2;
					out<=194;
				end
				if(in == 574) begin
					state<=2;
					out<=195;
				end
				if(in == 575) begin
					state<=2;
					out<=196;
				end
				if(in == 576) begin
					state<=2;
					out<=197;
				end
				if(in == 577) begin
					state<=2;
					out<=198;
				end
				if(in == 578) begin
					state<=2;
					out<=199;
				end
				if(in == 579) begin
					state<=2;
					out<=200;
				end
				if(in == 580) begin
					state<=2;
					out<=201;
				end
				if(in == 581) begin
					state<=3;
					out<=202;
				end
				if(in == 582) begin
					state<=5;
					out<=203;
				end
				if(in == 583) begin
					state<=3;
					out<=204;
				end
				if(in == 584) begin
					state<=5;
					out<=205;
				end
				if(in == 585) begin
					state<=3;
					out<=206;
				end
				if(in == 586) begin
					state<=5;
					out<=207;
				end
				if(in == 587) begin
					state<=5;
					out<=208;
				end
				if(in == 588) begin
					state<=5;
					out<=209;
				end
				if(in == 589) begin
					state<=5;
					out<=210;
				end
				if(in == 590) begin
					state<=5;
					out<=211;
				end
				if(in == 591) begin
					state<=5;
					out<=212;
				end
				if(in == 592) begin
					state<=5;
					out<=213;
				end
				if(in == 593) begin
					state<=5;
					out<=214;
				end
				if(in == 594) begin
					state<=5;
					out<=215;
				end
				if(in == 595) begin
					state<=5;
					out<=216;
				end
				if(in == 596) begin
					state<=5;
					out<=217;
				end
				if(in == 597) begin
					state<=5;
					out<=218;
				end
				if(in == 598) begin
					state<=5;
					out<=219;
				end
				if(in == 599) begin
					state<=5;
					out<=220;
				end
				if(in == 600) begin
					state<=5;
					out<=221;
				end
				if(in == 601) begin
					state<=6;
					out<=222;
				end
				if(in == 602) begin
					state<=6;
					out<=223;
				end
				if(in == 603) begin
					state<=6;
					out<=224;
				end
				if(in == 604) begin
					state<=6;
					out<=225;
				end
				if(in == 605) begin
					state<=6;
					out<=226;
				end
				if(in == 606) begin
					state<=6;
					out<=227;
				end
				if(in == 607) begin
					state<=6;
					out<=228;
				end
				if(in == 608) begin
					state<=6;
					out<=229;
				end
				if(in == 609) begin
					state<=6;
					out<=230;
				end
				if(in == 610) begin
					state<=6;
					out<=231;
				end
				if(in == 611) begin
					state<=6;
					out<=232;
				end
				if(in == 612) begin
					state<=6;
					out<=233;
				end
				if(in == 613) begin
					state<=6;
					out<=234;
				end
				if(in == 614) begin
					state<=6;
					out<=235;
				end
				if(in == 615) begin
					state<=6;
					out<=236;
				end
				if(in == 616) begin
					state<=6;
					out<=237;
				end
				if(in == 617) begin
					state<=5;
					out<=238;
				end
				if(in == 618) begin
					state<=5;
					out<=239;
				end
				if(in == 619) begin
					state<=5;
					out<=240;
				end
				if(in == 620) begin
					state<=5;
					out<=241;
				end
				if(in == 621) begin
					state<=5;
					out<=242;
				end
				if(in == 622) begin
					state<=5;
					out<=243;
				end
				if(in == 623) begin
					state<=5;
					out<=244;
				end
				if(in == 624) begin
					state<=5;
					out<=245;
				end
				if(in == 625) begin
					state<=5;
					out<=246;
				end
				if(in == 626) begin
					state<=5;
					out<=247;
				end
				if(in == 627) begin
					state<=5;
					out<=248;
				end
				if(in == 628) begin
					state<=5;
					out<=249;
				end
				if(in == 629) begin
					state<=5;
					out<=250;
				end
				if(in == 630) begin
					state<=5;
					out<=251;
				end
				if(in == 631) begin
					state<=5;
					out<=252;
				end
				if(in == 632) begin
					state<=5;
					out<=253;
				end
				if(in == 633) begin
					state<=3;
					out<=254;
				end
				if(in == 634) begin
					state<=5;
					out<=255;
				end
				if(in == 635) begin
					state<=3;
					out<=0;
				end
				if(in == 636) begin
					state<=5;
					out<=1;
				end
				if(in == 637) begin
					state<=3;
					out<=2;
				end
				if(in == 638) begin
					state<=5;
					out<=3;
				end
				if(in == 639) begin
					state<=5;
					out<=4;
				end
				if(in == 640) begin
					state<=5;
					out<=5;
				end
				if(in == 641) begin
					state<=5;
					out<=6;
				end
				if(in == 642) begin
					state<=5;
					out<=7;
				end
				if(in == 643) begin
					state<=5;
					out<=8;
				end
				if(in == 644) begin
					state<=5;
					out<=9;
				end
				if(in == 645) begin
					state<=5;
					out<=10;
				end
				if(in == 646) begin
					state<=5;
					out<=11;
				end
				if(in == 647) begin
					state<=5;
					out<=12;
				end
				if(in == 648) begin
					state<=5;
					out<=13;
				end
				if(in == 649) begin
					state<=5;
					out<=14;
				end
				if(in == 650) begin
					state<=5;
					out<=15;
				end
				if(in == 651) begin
					state<=5;
					out<=16;
				end
				if(in == 652) begin
					state<=5;
					out<=17;
				end
				if(in == 653) begin
					state<=6;
					out<=18;
				end
				if(in == 654) begin
					state<=6;
					out<=19;
				end
				if(in == 655) begin
					state<=6;
					out<=20;
				end
				if(in == 656) begin
					state<=6;
					out<=21;
				end
				if(in == 657) begin
					state<=6;
					out<=22;
				end
				if(in == 658) begin
					state<=6;
					out<=23;
				end
				if(in == 659) begin
					state<=6;
					out<=24;
				end
				if(in == 660) begin
					state<=6;
					out<=25;
				end
				if(in == 661) begin
					state<=6;
					out<=26;
				end
				if(in == 662) begin
					state<=6;
					out<=27;
				end
				if(in == 663) begin
					state<=6;
					out<=28;
				end
				if(in == 664) begin
					state<=6;
					out<=29;
				end
				if(in == 665) begin
					state<=6;
					out<=30;
				end
				if(in == 666) begin
					state<=6;
					out<=31;
				end
				if(in == 667) begin
					state<=6;
					out<=32;
				end
				if(in == 668) begin
					state<=6;
					out<=33;
				end
				if(in == 669) begin
					state<=5;
					out<=34;
				end
				if(in == 670) begin
					state<=5;
					out<=35;
				end
				if(in == 671) begin
					state<=5;
					out<=36;
				end
				if(in == 672) begin
					state<=5;
					out<=37;
				end
				if(in == 673) begin
					state<=5;
					out<=38;
				end
				if(in == 674) begin
					state<=5;
					out<=39;
				end
				if(in == 675) begin
					state<=5;
					out<=40;
				end
				if(in == 676) begin
					state<=5;
					out<=41;
				end
				if(in == 677) begin
					state<=5;
					out<=42;
				end
				if(in == 678) begin
					state<=5;
					out<=43;
				end
				if(in == 679) begin
					state<=5;
					out<=44;
				end
				if(in == 680) begin
					state<=5;
					out<=45;
				end
				if(in == 681) begin
					state<=5;
					out<=46;
				end
				if(in == 682) begin
					state<=5;
					out<=47;
				end
				if(in == 683) begin
					state<=5;
					out<=48;
				end
				if(in == 684) begin
					state<=5;
					out<=49;
				end
				if(in == 685) begin
					state<=2;
					out<=50;
				end
				if(in == 686) begin
					state<=2;
					out<=51;
				end
				if(in == 687) begin
					state<=2;
					out<=52;
				end
				if(in == 688) begin
					state<=2;
					out<=53;
				end
				if(in == 689) begin
					state<=2;
					out<=54;
				end
				if(in == 690) begin
					state<=2;
					out<=55;
				end
				if(in == 691) begin
					state<=2;
					out<=56;
				end
				if(in == 692) begin
					state<=2;
					out<=57;
				end
				if(in == 693) begin
					state<=2;
					out<=58;
				end
				if(in == 694) begin
					state<=2;
					out<=59;
				end
				if(in == 695) begin
					state<=2;
					out<=60;
				end
				if(in == 696) begin
					state<=2;
					out<=61;
				end
				if(in == 697) begin
					state<=3;
					out<=62;
				end
				if(in == 698) begin
					state<=5;
					out<=63;
				end
				if(in == 699) begin
					state<=3;
					out<=64;
				end
				if(in == 700) begin
					state<=5;
					out<=65;
				end
				if(in == 701) begin
					state<=3;
					out<=66;
				end
				if(in == 702) begin
					state<=5;
					out<=67;
				end
				if(in == 703) begin
					state<=5;
					out<=68;
				end
				if(in == 704) begin
					state<=5;
					out<=69;
				end
				if(in == 705) begin
					state<=5;
					out<=70;
				end
				if(in == 706) begin
					state<=5;
					out<=71;
				end
				if(in == 707) begin
					state<=5;
					out<=72;
				end
				if(in == 708) begin
					state<=5;
					out<=73;
				end
				if(in == 709) begin
					state<=5;
					out<=74;
				end
				if(in == 710) begin
					state<=5;
					out<=75;
				end
				if(in == 711) begin
					state<=5;
					out<=76;
				end
				if(in == 712) begin
					state<=5;
					out<=77;
				end
				if(in == 713) begin
					state<=5;
					out<=78;
				end
				if(in == 714) begin
					state<=5;
					out<=79;
				end
				if(in == 715) begin
					state<=5;
					out<=80;
				end
				if(in == 716) begin
					state<=5;
					out<=81;
				end
				if(in == 717) begin
					state<=6;
					out<=82;
				end
				if(in == 718) begin
					state<=6;
					out<=83;
				end
				if(in == 719) begin
					state<=6;
					out<=84;
				end
				if(in == 720) begin
					state<=6;
					out<=85;
				end
				if(in == 721) begin
					state<=6;
					out<=86;
				end
				if(in == 722) begin
					state<=6;
					out<=87;
				end
				if(in == 723) begin
					state<=6;
					out<=88;
				end
				if(in == 724) begin
					state<=6;
					out<=89;
				end
				if(in == 725) begin
					state<=6;
					out<=90;
				end
				if(in == 726) begin
					state<=6;
					out<=91;
				end
				if(in == 727) begin
					state<=6;
					out<=92;
				end
				if(in == 728) begin
					state<=6;
					out<=93;
				end
				if(in == 729) begin
					state<=6;
					out<=94;
				end
				if(in == 730) begin
					state<=6;
					out<=95;
				end
				if(in == 731) begin
					state<=6;
					out<=96;
				end
				if(in == 732) begin
					state<=6;
					out<=97;
				end
				if(in == 733) begin
					state<=5;
					out<=98;
				end
				if(in == 734) begin
					state<=5;
					out<=99;
				end
				if(in == 735) begin
					state<=5;
					out<=100;
				end
				if(in == 736) begin
					state<=5;
					out<=101;
				end
				if(in == 737) begin
					state<=5;
					out<=102;
				end
				if(in == 738) begin
					state<=5;
					out<=103;
				end
				if(in == 739) begin
					state<=5;
					out<=104;
				end
				if(in == 740) begin
					state<=5;
					out<=105;
				end
				if(in == 741) begin
					state<=5;
					out<=106;
				end
				if(in == 742) begin
					state<=5;
					out<=107;
				end
				if(in == 743) begin
					state<=5;
					out<=108;
				end
				if(in == 744) begin
					state<=5;
					out<=109;
				end
				if(in == 745) begin
					state<=5;
					out<=110;
				end
				if(in == 746) begin
					state<=5;
					out<=111;
				end
				if(in == 747) begin
					state<=5;
					out<=112;
				end
				if(in == 748) begin
					state<=5;
					out<=113;
				end
				if(in == 749) begin
					state<=3;
					out<=114;
				end
				if(in == 750) begin
					state<=5;
					out<=115;
				end
				if(in == 751) begin
					state<=3;
					out<=116;
				end
				if(in == 752) begin
					state<=5;
					out<=117;
				end
				if(in == 753) begin
					state<=3;
					out<=118;
				end
				if(in == 754) begin
					state<=5;
					out<=119;
				end
				if(in == 755) begin
					state<=5;
					out<=120;
				end
				if(in == 756) begin
					state<=5;
					out<=121;
				end
				if(in == 757) begin
					state<=5;
					out<=122;
				end
				if(in == 758) begin
					state<=5;
					out<=123;
				end
				if(in == 759) begin
					state<=5;
					out<=124;
				end
				if(in == 760) begin
					state<=5;
					out<=125;
				end
				if(in == 761) begin
					state<=5;
					out<=126;
				end
				if(in == 762) begin
					state<=5;
					out<=127;
				end
				if(in == 763) begin
					state<=5;
					out<=128;
				end
				if(in == 764) begin
					state<=5;
					out<=129;
				end
				if(in == 765) begin
					state<=5;
					out<=130;
				end
				if(in == 766) begin
					state<=5;
					out<=131;
				end
				if(in == 767) begin
					state<=5;
					out<=132;
				end
				if(in == 768) begin
					state<=5;
					out<=133;
				end
				if(in == 769) begin
					state<=6;
					out<=134;
				end
				if(in == 770) begin
					state<=6;
					out<=135;
				end
				if(in == 771) begin
					state<=6;
					out<=136;
				end
				if(in == 772) begin
					state<=6;
					out<=137;
				end
				if(in == 773) begin
					state<=6;
					out<=138;
				end
				if(in == 774) begin
					state<=6;
					out<=139;
				end
				if(in == 775) begin
					state<=6;
					out<=140;
				end
				if(in == 776) begin
					state<=6;
					out<=141;
				end
				if(in == 777) begin
					state<=6;
					out<=142;
				end
				if(in == 778) begin
					state<=6;
					out<=143;
				end
				if(in == 779) begin
					state<=6;
					out<=144;
				end
				if(in == 780) begin
					state<=6;
					out<=145;
				end
				if(in == 781) begin
					state<=6;
					out<=146;
				end
				if(in == 782) begin
					state<=6;
					out<=147;
				end
				if(in == 783) begin
					state<=6;
					out<=148;
				end
				if(in == 784) begin
					state<=6;
					out<=149;
				end
				if(in == 785) begin
					state<=5;
					out<=150;
				end
				if(in == 786) begin
					state<=5;
					out<=151;
				end
				if(in == 787) begin
					state<=5;
					out<=152;
				end
				if(in == 788) begin
					state<=5;
					out<=153;
				end
				if(in == 789) begin
					state<=5;
					out<=154;
				end
				if(in == 790) begin
					state<=5;
					out<=155;
				end
				if(in == 791) begin
					state<=5;
					out<=156;
				end
				if(in == 792) begin
					state<=5;
					out<=157;
				end
				if(in == 793) begin
					state<=5;
					out<=158;
				end
				if(in == 794) begin
					state<=5;
					out<=159;
				end
				if(in == 795) begin
					state<=5;
					out<=160;
				end
				if(in == 796) begin
					state<=5;
					out<=161;
				end
				if(in == 797) begin
					state<=5;
					out<=162;
				end
				if(in == 798) begin
					state<=5;
					out<=163;
				end
				if(in == 799) begin
					state<=5;
					out<=164;
				end
				if(in == 800) begin
					state<=5;
					out<=165;
				end
				if(in == 801) begin
					state<=2;
					out<=166;
				end
				if(in == 802) begin
					state<=2;
					out<=167;
				end
				if(in == 803) begin
					state<=2;
					out<=168;
				end
				if(in == 804) begin
					state<=2;
					out<=169;
				end
				if(in == 805) begin
					state<=2;
					out<=170;
				end
				if(in == 806) begin
					state<=2;
					out<=171;
				end
				if(in == 807) begin
					state<=2;
					out<=172;
				end
				if(in == 808) begin
					state<=2;
					out<=173;
				end
				if(in == 809) begin
					state<=2;
					out<=174;
				end
				if(in == 810) begin
					state<=2;
					out<=175;
				end
				if(in == 811) begin
					state<=2;
					out<=176;
				end
				if(in == 812) begin
					state<=2;
					out<=177;
				end
				if(in == 813) begin
					state<=3;
					out<=178;
				end
				if(in == 814) begin
					state<=5;
					out<=179;
				end
				if(in == 815) begin
					state<=3;
					out<=180;
				end
				if(in == 816) begin
					state<=5;
					out<=181;
				end
				if(in == 817) begin
					state<=3;
					out<=182;
				end
				if(in == 818) begin
					state<=5;
					out<=183;
				end
				if(in == 819) begin
					state<=5;
					out<=184;
				end
				if(in == 820) begin
					state<=5;
					out<=185;
				end
				if(in == 821) begin
					state<=5;
					out<=186;
				end
				if(in == 822) begin
					state<=5;
					out<=187;
				end
				if(in == 823) begin
					state<=5;
					out<=188;
				end
				if(in == 824) begin
					state<=5;
					out<=189;
				end
				if(in == 825) begin
					state<=5;
					out<=190;
				end
				if(in == 826) begin
					state<=5;
					out<=191;
				end
				if(in == 827) begin
					state<=5;
					out<=192;
				end
				if(in == 828) begin
					state<=5;
					out<=193;
				end
				if(in == 829) begin
					state<=5;
					out<=194;
				end
				if(in == 830) begin
					state<=5;
					out<=195;
				end
				if(in == 831) begin
					state<=5;
					out<=196;
				end
				if(in == 832) begin
					state<=5;
					out<=197;
				end
				if(in == 833) begin
					state<=6;
					out<=198;
				end
				if(in == 834) begin
					state<=6;
					out<=199;
				end
				if(in == 835) begin
					state<=6;
					out<=200;
				end
				if(in == 836) begin
					state<=6;
					out<=201;
				end
				if(in == 837) begin
					state<=6;
					out<=202;
				end
				if(in == 838) begin
					state<=6;
					out<=203;
				end
				if(in == 839) begin
					state<=6;
					out<=204;
				end
				if(in == 840) begin
					state<=6;
					out<=205;
				end
				if(in == 841) begin
					state<=6;
					out<=206;
				end
				if(in == 842) begin
					state<=6;
					out<=207;
				end
				if(in == 843) begin
					state<=6;
					out<=208;
				end
				if(in == 844) begin
					state<=6;
					out<=209;
				end
				if(in == 845) begin
					state<=6;
					out<=210;
				end
				if(in == 846) begin
					state<=6;
					out<=211;
				end
				if(in == 847) begin
					state<=6;
					out<=212;
				end
				if(in == 848) begin
					state<=6;
					out<=213;
				end
				if(in == 849) begin
					state<=5;
					out<=214;
				end
				if(in == 850) begin
					state<=5;
					out<=215;
				end
				if(in == 851) begin
					state<=5;
					out<=216;
				end
				if(in == 852) begin
					state<=5;
					out<=217;
				end
				if(in == 853) begin
					state<=5;
					out<=218;
				end
				if(in == 854) begin
					state<=5;
					out<=219;
				end
				if(in == 855) begin
					state<=5;
					out<=220;
				end
				if(in == 856) begin
					state<=5;
					out<=221;
				end
				if(in == 857) begin
					state<=5;
					out<=222;
				end
				if(in == 858) begin
					state<=5;
					out<=223;
				end
				if(in == 859) begin
					state<=5;
					out<=224;
				end
				if(in == 860) begin
					state<=5;
					out<=225;
				end
				if(in == 861) begin
					state<=5;
					out<=226;
				end
				if(in == 862) begin
					state<=5;
					out<=227;
				end
				if(in == 863) begin
					state<=5;
					out<=228;
				end
				if(in == 864) begin
					state<=5;
					out<=229;
				end
				if(in == 865) begin
					state<=3;
					out<=230;
				end
				if(in == 866) begin
					state<=5;
					out<=231;
				end
				if(in == 867) begin
					state<=3;
					out<=232;
				end
				if(in == 868) begin
					state<=5;
					out<=233;
				end
				if(in == 869) begin
					state<=3;
					out<=234;
				end
				if(in == 870) begin
					state<=5;
					out<=235;
				end
				if(in == 871) begin
					state<=5;
					out<=236;
				end
				if(in == 872) begin
					state<=5;
					out<=237;
				end
				if(in == 873) begin
					state<=5;
					out<=238;
				end
				if(in == 874) begin
					state<=5;
					out<=239;
				end
				if(in == 875) begin
					state<=5;
					out<=240;
				end
				if(in == 876) begin
					state<=5;
					out<=241;
				end
				if(in == 877) begin
					state<=5;
					out<=242;
				end
				if(in == 878) begin
					state<=5;
					out<=243;
				end
				if(in == 879) begin
					state<=5;
					out<=244;
				end
				if(in == 880) begin
					state<=5;
					out<=245;
				end
				if(in == 881) begin
					state<=5;
					out<=246;
				end
				if(in == 882) begin
					state<=5;
					out<=247;
				end
				if(in == 883) begin
					state<=5;
					out<=248;
				end
				if(in == 884) begin
					state<=5;
					out<=249;
				end
				if(in == 885) begin
					state<=6;
					out<=250;
				end
				if(in == 886) begin
					state<=6;
					out<=251;
				end
				if(in == 887) begin
					state<=6;
					out<=252;
				end
				if(in == 888) begin
					state<=6;
					out<=253;
				end
				if(in == 889) begin
					state<=6;
					out<=254;
				end
				if(in == 890) begin
					state<=6;
					out<=255;
				end
				if(in == 891) begin
					state<=6;
					out<=0;
				end
				if(in == 892) begin
					state<=6;
					out<=1;
				end
				if(in == 893) begin
					state<=6;
					out<=2;
				end
				if(in == 894) begin
					state<=6;
					out<=3;
				end
				if(in == 895) begin
					state<=6;
					out<=4;
				end
				if(in == 896) begin
					state<=6;
					out<=5;
				end
				if(in == 897) begin
					state<=6;
					out<=6;
				end
				if(in == 898) begin
					state<=6;
					out<=7;
				end
				if(in == 899) begin
					state<=6;
					out<=8;
				end
				if(in == 900) begin
					state<=6;
					out<=9;
				end
				if(in == 901) begin
					state<=5;
					out<=10;
				end
				if(in == 902) begin
					state<=5;
					out<=11;
				end
				if(in == 903) begin
					state<=5;
					out<=12;
				end
				if(in == 904) begin
					state<=5;
					out<=13;
				end
				if(in == 905) begin
					state<=5;
					out<=14;
				end
				if(in == 906) begin
					state<=5;
					out<=15;
				end
				if(in == 907) begin
					state<=5;
					out<=16;
				end
				if(in == 908) begin
					state<=5;
					out<=17;
				end
				if(in == 909) begin
					state<=5;
					out<=18;
				end
				if(in == 910) begin
					state<=5;
					out<=19;
				end
				if(in == 911) begin
					state<=5;
					out<=20;
				end
				if(in == 912) begin
					state<=5;
					out<=21;
				end
				if(in == 913) begin
					state<=5;
					out<=22;
				end
				if(in == 914) begin
					state<=5;
					out<=23;
				end
				if(in == 915) begin
					state<=5;
					out<=24;
				end
				if(in == 916) begin
					state<=5;
					out<=25;
				end
				if(in == 917) begin
					state<=2;
					out<=26;
				end
				if(in == 918) begin
					state<=2;
					out<=27;
				end
				if(in == 919) begin
					state<=2;
					out<=28;
				end
				if(in == 920) begin
					state<=2;
					out<=29;
				end
				if(in == 921) begin
					state<=2;
					out<=30;
				end
				if(in == 922) begin
					state<=2;
					out<=31;
				end
				if(in == 923) begin
					state<=2;
					out<=32;
				end
				if(in == 924) begin
					state<=2;
					out<=33;
				end
				if(in == 925) begin
					state<=2;
					out<=34;
				end
				if(in == 926) begin
					state<=2;
					out<=35;
				end
				if(in == 927) begin
					state<=2;
					out<=36;
				end
				if(in == 928) begin
					state<=2;
					out<=37;
				end
			end
			6: begin
				if(in == 0) begin
					state<=3;
					out<=38;
				end
				if(in == 1) begin
					state<=1;
					out<=39;
				end
				if(in == 2) begin
					state<=6;
					out<=40;
				end
				if(in == 3) begin
					state<=3;
					out<=41;
				end
				if(in == 4) begin
					state<=7;
					out<=42;
				end
				if(in == 5) begin
					state<=3;
					out<=43;
				end
				if(in == 6) begin
					state<=7;
					out<=44;
				end
				if(in == 7) begin
					state<=7;
					out<=45;
				end
				if(in == 8) begin
					state<=7;
					out<=46;
				end
				if(in == 9) begin
					state<=7;
					out<=47;
				end
				if(in == 10) begin
					state<=7;
					out<=48;
				end
				if(in == 11) begin
					state<=7;
					out<=49;
				end
				if(in == 12) begin
					state<=7;
					out<=50;
				end
				if(in == 13) begin
					state<=7;
					out<=51;
				end
				if(in == 14) begin
					state<=7;
					out<=52;
				end
				if(in == 15) begin
					state<=7;
					out<=53;
				end
				if(in == 16) begin
					state<=7;
					out<=54;
				end
				if(in == 17) begin
					state<=7;
					out<=55;
				end
				if(in == 18) begin
					state<=7;
					out<=56;
				end
				if(in == 19) begin
					state<=7;
					out<=57;
				end
				if(in == 20) begin
					state<=7;
					out<=58;
				end
				if(in == 21) begin
					state<=7;
					out<=59;
				end
				if(in == 22) begin
					state<=7;
					out<=60;
				end
				if(in == 23) begin
					state<=7;
					out<=61;
				end
				if(in == 24) begin
					state<=7;
					out<=62;
				end
				if(in == 25) begin
					state<=7;
					out<=63;
				end
				if(in == 26) begin
					state<=7;
					out<=64;
				end
				if(in == 27) begin
					state<=7;
					out<=65;
				end
				if(in == 28) begin
					state<=7;
					out<=66;
				end
				if(in == 29) begin
					state<=7;
					out<=67;
				end
				if(in == 30) begin
					state<=7;
					out<=68;
				end
				if(in == 31) begin
					state<=7;
					out<=69;
				end
				if(in == 32) begin
					state<=7;
					out<=70;
				end
				if(in == 33) begin
					state<=7;
					out<=71;
				end
				if(in == 34) begin
					state<=7;
					out<=72;
				end
				if(in == 35) begin
					state<=7;
					out<=73;
				end
				if(in == 36) begin
					state<=7;
					out<=74;
				end
				if(in == 37) begin
					state<=7;
					out<=75;
				end
				if(in == 38) begin
					state<=7;
					out<=76;
				end
				if(in == 39) begin
					state<=7;
					out<=77;
				end
				if(in == 40) begin
					state<=7;
					out<=78;
				end
				if(in == 41) begin
					state<=7;
					out<=79;
				end
				if(in == 42) begin
					state<=7;
					out<=80;
				end
				if(in == 43) begin
					state<=7;
					out<=81;
				end
				if(in == 44) begin
					state<=7;
					out<=82;
				end
				if(in == 45) begin
					state<=7;
					out<=83;
				end
				if(in == 46) begin
					state<=7;
					out<=84;
				end
				if(in == 47) begin
					state<=7;
					out<=85;
				end
				if(in == 48) begin
					state<=7;
					out<=86;
				end
				if(in == 49) begin
					state<=7;
					out<=87;
				end
				if(in == 50) begin
					state<=7;
					out<=88;
				end
				if(in == 51) begin
					state<=7;
					out<=89;
				end
				if(in == 52) begin
					state<=7;
					out<=90;
				end
				if(in == 53) begin
					state<=3;
					out<=91;
				end
				if(in == 54) begin
					state<=6;
					out<=92;
				end
				if(in == 55) begin
					state<=3;
					out<=93;
				end
				if(in == 56) begin
					state<=7;
					out<=94;
				end
				if(in == 57) begin
					state<=3;
					out<=95;
				end
				if(in == 58) begin
					state<=7;
					out<=96;
				end
				if(in == 59) begin
					state<=7;
					out<=97;
				end
				if(in == 60) begin
					state<=7;
					out<=98;
				end
				if(in == 61) begin
					state<=7;
					out<=99;
				end
				if(in == 62) begin
					state<=7;
					out<=100;
				end
				if(in == 63) begin
					state<=7;
					out<=101;
				end
				if(in == 64) begin
					state<=7;
					out<=102;
				end
				if(in == 65) begin
					state<=7;
					out<=103;
				end
				if(in == 66) begin
					state<=7;
					out<=104;
				end
				if(in == 67) begin
					state<=7;
					out<=105;
				end
				if(in == 68) begin
					state<=7;
					out<=106;
				end
				if(in == 69) begin
					state<=7;
					out<=107;
				end
				if(in == 70) begin
					state<=7;
					out<=108;
				end
				if(in == 71) begin
					state<=7;
					out<=109;
				end
				if(in == 72) begin
					state<=7;
					out<=110;
				end
				if(in == 73) begin
					state<=7;
					out<=111;
				end
				if(in == 74) begin
					state<=7;
					out<=112;
				end
				if(in == 75) begin
					state<=7;
					out<=113;
				end
				if(in == 76) begin
					state<=7;
					out<=114;
				end
				if(in == 77) begin
					state<=7;
					out<=115;
				end
				if(in == 78) begin
					state<=7;
					out<=116;
				end
				if(in == 79) begin
					state<=7;
					out<=117;
				end
				if(in == 80) begin
					state<=7;
					out<=118;
				end
				if(in == 81) begin
					state<=7;
					out<=119;
				end
				if(in == 82) begin
					state<=7;
					out<=120;
				end
				if(in == 83) begin
					state<=7;
					out<=121;
				end
				if(in == 84) begin
					state<=7;
					out<=122;
				end
				if(in == 85) begin
					state<=7;
					out<=123;
				end
				if(in == 86) begin
					state<=7;
					out<=124;
				end
				if(in == 87) begin
					state<=7;
					out<=125;
				end
				if(in == 88) begin
					state<=7;
					out<=126;
				end
				if(in == 89) begin
					state<=7;
					out<=127;
				end
				if(in == 90) begin
					state<=7;
					out<=128;
				end
				if(in == 91) begin
					state<=7;
					out<=129;
				end
				if(in == 92) begin
					state<=7;
					out<=130;
				end
				if(in == 93) begin
					state<=7;
					out<=131;
				end
				if(in == 94) begin
					state<=7;
					out<=132;
				end
				if(in == 95) begin
					state<=7;
					out<=133;
				end
				if(in == 96) begin
					state<=7;
					out<=134;
				end
				if(in == 97) begin
					state<=7;
					out<=135;
				end
				if(in == 98) begin
					state<=7;
					out<=136;
				end
				if(in == 99) begin
					state<=7;
					out<=137;
				end
				if(in == 100) begin
					state<=7;
					out<=138;
				end
				if(in == 101) begin
					state<=7;
					out<=139;
				end
				if(in == 102) begin
					state<=7;
					out<=140;
				end
				if(in == 103) begin
					state<=7;
					out<=141;
				end
				if(in == 104) begin
					state<=7;
					out<=142;
				end
				if(in == 105) begin
					state<=2;
					out<=143;
				end
				if(in == 106) begin
					state<=2;
					out<=144;
				end
				if(in == 107) begin
					state<=2;
					out<=145;
				end
				if(in == 108) begin
					state<=2;
					out<=146;
				end
				if(in == 109) begin
					state<=2;
					out<=147;
				end
				if(in == 110) begin
					state<=2;
					out<=148;
				end
				if(in == 111) begin
					state<=2;
					out<=149;
				end
				if(in == 112) begin
					state<=2;
					out<=150;
				end
				if(in == 113) begin
					state<=2;
					out<=151;
				end
				if(in == 114) begin
					state<=2;
					out<=152;
				end
				if(in == 115) begin
					state<=2;
					out<=153;
				end
				if(in == 116) begin
					state<=2;
					out<=154;
				end
				if(in == 117) begin
					state<=3;
					out<=155;
				end
				if(in == 118) begin
					state<=6;
					out<=156;
				end
				if(in == 119) begin
					state<=3;
					out<=157;
				end
				if(in == 120) begin
					state<=7;
					out<=158;
				end
				if(in == 121) begin
					state<=3;
					out<=159;
				end
				if(in == 122) begin
					state<=7;
					out<=160;
				end
				if(in == 123) begin
					state<=7;
					out<=161;
				end
				if(in == 124) begin
					state<=7;
					out<=162;
				end
				if(in == 125) begin
					state<=7;
					out<=163;
				end
				if(in == 126) begin
					state<=7;
					out<=164;
				end
				if(in == 127) begin
					state<=7;
					out<=165;
				end
				if(in == 128) begin
					state<=7;
					out<=166;
				end
				if(in == 129) begin
					state<=7;
					out<=167;
				end
				if(in == 130) begin
					state<=7;
					out<=168;
				end
				if(in == 131) begin
					state<=7;
					out<=169;
				end
				if(in == 132) begin
					state<=7;
					out<=170;
				end
				if(in == 133) begin
					state<=7;
					out<=171;
				end
				if(in == 134) begin
					state<=7;
					out<=172;
				end
				if(in == 135) begin
					state<=7;
					out<=173;
				end
				if(in == 136) begin
					state<=7;
					out<=174;
				end
				if(in == 137) begin
					state<=7;
					out<=175;
				end
				if(in == 138) begin
					state<=7;
					out<=176;
				end
				if(in == 139) begin
					state<=7;
					out<=177;
				end
				if(in == 140) begin
					state<=7;
					out<=178;
				end
				if(in == 141) begin
					state<=7;
					out<=179;
				end
				if(in == 142) begin
					state<=7;
					out<=180;
				end
				if(in == 143) begin
					state<=7;
					out<=181;
				end
				if(in == 144) begin
					state<=7;
					out<=182;
				end
				if(in == 145) begin
					state<=7;
					out<=183;
				end
				if(in == 146) begin
					state<=7;
					out<=184;
				end
				if(in == 147) begin
					state<=7;
					out<=185;
				end
				if(in == 148) begin
					state<=7;
					out<=186;
				end
				if(in == 149) begin
					state<=7;
					out<=187;
				end
				if(in == 150) begin
					state<=7;
					out<=188;
				end
				if(in == 151) begin
					state<=7;
					out<=189;
				end
				if(in == 152) begin
					state<=7;
					out<=190;
				end
				if(in == 153) begin
					state<=7;
					out<=191;
				end
				if(in == 154) begin
					state<=7;
					out<=192;
				end
				if(in == 155) begin
					state<=7;
					out<=193;
				end
				if(in == 156) begin
					state<=7;
					out<=194;
				end
				if(in == 157) begin
					state<=7;
					out<=195;
				end
				if(in == 158) begin
					state<=7;
					out<=196;
				end
				if(in == 159) begin
					state<=7;
					out<=197;
				end
				if(in == 160) begin
					state<=7;
					out<=198;
				end
				if(in == 161) begin
					state<=7;
					out<=199;
				end
				if(in == 162) begin
					state<=7;
					out<=200;
				end
				if(in == 163) begin
					state<=7;
					out<=201;
				end
				if(in == 164) begin
					state<=7;
					out<=202;
				end
				if(in == 165) begin
					state<=7;
					out<=203;
				end
				if(in == 166) begin
					state<=7;
					out<=204;
				end
				if(in == 167) begin
					state<=7;
					out<=205;
				end
				if(in == 168) begin
					state<=7;
					out<=206;
				end
				if(in == 169) begin
					state<=3;
					out<=207;
				end
				if(in == 170) begin
					state<=6;
					out<=208;
				end
				if(in == 171) begin
					state<=3;
					out<=209;
				end
				if(in == 172) begin
					state<=7;
					out<=210;
				end
				if(in == 173) begin
					state<=3;
					out<=211;
				end
				if(in == 174) begin
					state<=7;
					out<=212;
				end
				if(in == 175) begin
					state<=7;
					out<=213;
				end
				if(in == 176) begin
					state<=7;
					out<=214;
				end
				if(in == 177) begin
					state<=7;
					out<=215;
				end
				if(in == 178) begin
					state<=7;
					out<=216;
				end
				if(in == 179) begin
					state<=7;
					out<=217;
				end
				if(in == 180) begin
					state<=7;
					out<=218;
				end
				if(in == 181) begin
					state<=7;
					out<=219;
				end
				if(in == 182) begin
					state<=7;
					out<=220;
				end
				if(in == 183) begin
					state<=7;
					out<=221;
				end
				if(in == 184) begin
					state<=7;
					out<=222;
				end
				if(in == 185) begin
					state<=7;
					out<=223;
				end
				if(in == 186) begin
					state<=7;
					out<=224;
				end
				if(in == 187) begin
					state<=7;
					out<=225;
				end
				if(in == 188) begin
					state<=7;
					out<=226;
				end
				if(in == 189) begin
					state<=7;
					out<=227;
				end
				if(in == 190) begin
					state<=7;
					out<=228;
				end
				if(in == 191) begin
					state<=7;
					out<=229;
				end
				if(in == 192) begin
					state<=7;
					out<=230;
				end
				if(in == 193) begin
					state<=7;
					out<=231;
				end
				if(in == 194) begin
					state<=7;
					out<=232;
				end
				if(in == 195) begin
					state<=7;
					out<=233;
				end
				if(in == 196) begin
					state<=7;
					out<=234;
				end
				if(in == 197) begin
					state<=7;
					out<=235;
				end
				if(in == 198) begin
					state<=7;
					out<=236;
				end
				if(in == 199) begin
					state<=7;
					out<=237;
				end
				if(in == 200) begin
					state<=7;
					out<=238;
				end
				if(in == 201) begin
					state<=7;
					out<=239;
				end
				if(in == 202) begin
					state<=7;
					out<=240;
				end
				if(in == 203) begin
					state<=7;
					out<=241;
				end
				if(in == 204) begin
					state<=7;
					out<=242;
				end
				if(in == 205) begin
					state<=7;
					out<=243;
				end
				if(in == 206) begin
					state<=7;
					out<=244;
				end
				if(in == 207) begin
					state<=7;
					out<=245;
				end
				if(in == 208) begin
					state<=7;
					out<=246;
				end
				if(in == 209) begin
					state<=7;
					out<=247;
				end
				if(in == 210) begin
					state<=7;
					out<=248;
				end
				if(in == 211) begin
					state<=7;
					out<=249;
				end
				if(in == 212) begin
					state<=7;
					out<=250;
				end
				if(in == 213) begin
					state<=7;
					out<=251;
				end
				if(in == 214) begin
					state<=7;
					out<=252;
				end
				if(in == 215) begin
					state<=7;
					out<=253;
				end
				if(in == 216) begin
					state<=7;
					out<=254;
				end
				if(in == 217) begin
					state<=7;
					out<=255;
				end
				if(in == 218) begin
					state<=7;
					out<=0;
				end
				if(in == 219) begin
					state<=7;
					out<=1;
				end
				if(in == 220) begin
					state<=7;
					out<=2;
				end
				if(in == 221) begin
					state<=2;
					out<=3;
				end
				if(in == 222) begin
					state<=2;
					out<=4;
				end
				if(in == 223) begin
					state<=2;
					out<=5;
				end
				if(in == 224) begin
					state<=2;
					out<=6;
				end
				if(in == 225) begin
					state<=2;
					out<=7;
				end
				if(in == 226) begin
					state<=2;
					out<=8;
				end
				if(in == 227) begin
					state<=2;
					out<=9;
				end
				if(in == 228) begin
					state<=2;
					out<=10;
				end
				if(in == 229) begin
					state<=2;
					out<=11;
				end
				if(in == 230) begin
					state<=2;
					out<=12;
				end
				if(in == 231) begin
					state<=2;
					out<=13;
				end
				if(in == 232) begin
					state<=2;
					out<=14;
				end
				if(in == 233) begin
					state<=3;
					out<=15;
				end
				if(in == 234) begin
					state<=6;
					out<=16;
				end
				if(in == 235) begin
					state<=3;
					out<=17;
				end
				if(in == 236) begin
					state<=7;
					out<=18;
				end
				if(in == 237) begin
					state<=3;
					out<=19;
				end
				if(in == 238) begin
					state<=7;
					out<=20;
				end
				if(in == 239) begin
					state<=7;
					out<=21;
				end
				if(in == 240) begin
					state<=7;
					out<=22;
				end
				if(in == 241) begin
					state<=7;
					out<=23;
				end
				if(in == 242) begin
					state<=7;
					out<=24;
				end
				if(in == 243) begin
					state<=7;
					out<=25;
				end
				if(in == 244) begin
					state<=7;
					out<=26;
				end
				if(in == 245) begin
					state<=7;
					out<=27;
				end
				if(in == 246) begin
					state<=7;
					out<=28;
				end
				if(in == 247) begin
					state<=7;
					out<=29;
				end
				if(in == 248) begin
					state<=7;
					out<=30;
				end
				if(in == 249) begin
					state<=7;
					out<=31;
				end
				if(in == 250) begin
					state<=7;
					out<=32;
				end
				if(in == 251) begin
					state<=7;
					out<=33;
				end
				if(in == 252) begin
					state<=7;
					out<=34;
				end
				if(in == 253) begin
					state<=7;
					out<=35;
				end
				if(in == 254) begin
					state<=7;
					out<=36;
				end
				if(in == 255) begin
					state<=7;
					out<=37;
				end
				if(in == 256) begin
					state<=7;
					out<=38;
				end
				if(in == 257) begin
					state<=7;
					out<=39;
				end
				if(in == 258) begin
					state<=7;
					out<=40;
				end
				if(in == 259) begin
					state<=7;
					out<=41;
				end
				if(in == 260) begin
					state<=7;
					out<=42;
				end
				if(in == 261) begin
					state<=7;
					out<=43;
				end
				if(in == 262) begin
					state<=7;
					out<=44;
				end
				if(in == 263) begin
					state<=7;
					out<=45;
				end
				if(in == 264) begin
					state<=7;
					out<=46;
				end
				if(in == 265) begin
					state<=7;
					out<=47;
				end
				if(in == 266) begin
					state<=7;
					out<=48;
				end
				if(in == 267) begin
					state<=7;
					out<=49;
				end
				if(in == 268) begin
					state<=7;
					out<=50;
				end
				if(in == 269) begin
					state<=7;
					out<=51;
				end
				if(in == 270) begin
					state<=7;
					out<=52;
				end
				if(in == 271) begin
					state<=7;
					out<=53;
				end
				if(in == 272) begin
					state<=7;
					out<=54;
				end
				if(in == 273) begin
					state<=7;
					out<=55;
				end
				if(in == 274) begin
					state<=7;
					out<=56;
				end
				if(in == 275) begin
					state<=7;
					out<=57;
				end
				if(in == 276) begin
					state<=7;
					out<=58;
				end
				if(in == 277) begin
					state<=7;
					out<=59;
				end
				if(in == 278) begin
					state<=7;
					out<=60;
				end
				if(in == 279) begin
					state<=7;
					out<=61;
				end
				if(in == 280) begin
					state<=7;
					out<=62;
				end
				if(in == 281) begin
					state<=7;
					out<=63;
				end
				if(in == 282) begin
					state<=7;
					out<=64;
				end
				if(in == 283) begin
					state<=7;
					out<=65;
				end
				if(in == 284) begin
					state<=7;
					out<=66;
				end
				if(in == 285) begin
					state<=3;
					out<=67;
				end
				if(in == 286) begin
					state<=6;
					out<=68;
				end
				if(in == 287) begin
					state<=3;
					out<=69;
				end
				if(in == 288) begin
					state<=7;
					out<=70;
				end
				if(in == 289) begin
					state<=3;
					out<=71;
				end
				if(in == 290) begin
					state<=7;
					out<=72;
				end
				if(in == 291) begin
					state<=7;
					out<=73;
				end
				if(in == 292) begin
					state<=7;
					out<=74;
				end
				if(in == 293) begin
					state<=7;
					out<=75;
				end
				if(in == 294) begin
					state<=7;
					out<=76;
				end
				if(in == 295) begin
					state<=7;
					out<=77;
				end
				if(in == 296) begin
					state<=7;
					out<=78;
				end
				if(in == 297) begin
					state<=7;
					out<=79;
				end
				if(in == 298) begin
					state<=7;
					out<=80;
				end
				if(in == 299) begin
					state<=7;
					out<=81;
				end
				if(in == 300) begin
					state<=7;
					out<=82;
				end
				if(in == 301) begin
					state<=7;
					out<=83;
				end
				if(in == 302) begin
					state<=7;
					out<=84;
				end
				if(in == 303) begin
					state<=7;
					out<=85;
				end
				if(in == 304) begin
					state<=7;
					out<=86;
				end
				if(in == 305) begin
					state<=7;
					out<=87;
				end
				if(in == 306) begin
					state<=7;
					out<=88;
				end
				if(in == 307) begin
					state<=7;
					out<=89;
				end
				if(in == 308) begin
					state<=7;
					out<=90;
				end
				if(in == 309) begin
					state<=7;
					out<=91;
				end
				if(in == 310) begin
					state<=7;
					out<=92;
				end
				if(in == 311) begin
					state<=7;
					out<=93;
				end
				if(in == 312) begin
					state<=7;
					out<=94;
				end
				if(in == 313) begin
					state<=7;
					out<=95;
				end
				if(in == 314) begin
					state<=7;
					out<=96;
				end
				if(in == 315) begin
					state<=7;
					out<=97;
				end
				if(in == 316) begin
					state<=7;
					out<=98;
				end
				if(in == 317) begin
					state<=7;
					out<=99;
				end
				if(in == 318) begin
					state<=7;
					out<=100;
				end
				if(in == 319) begin
					state<=7;
					out<=101;
				end
				if(in == 320) begin
					state<=7;
					out<=102;
				end
				if(in == 321) begin
					state<=7;
					out<=103;
				end
				if(in == 322) begin
					state<=7;
					out<=104;
				end
				if(in == 323) begin
					state<=7;
					out<=105;
				end
				if(in == 324) begin
					state<=7;
					out<=106;
				end
				if(in == 325) begin
					state<=7;
					out<=107;
				end
				if(in == 326) begin
					state<=7;
					out<=108;
				end
				if(in == 327) begin
					state<=7;
					out<=109;
				end
				if(in == 328) begin
					state<=7;
					out<=110;
				end
				if(in == 329) begin
					state<=7;
					out<=111;
				end
				if(in == 330) begin
					state<=7;
					out<=112;
				end
				if(in == 331) begin
					state<=7;
					out<=113;
				end
				if(in == 332) begin
					state<=7;
					out<=114;
				end
				if(in == 333) begin
					state<=7;
					out<=115;
				end
				if(in == 334) begin
					state<=7;
					out<=116;
				end
				if(in == 335) begin
					state<=7;
					out<=117;
				end
				if(in == 336) begin
					state<=7;
					out<=118;
				end
				if(in == 337) begin
					state<=2;
					out<=119;
				end
				if(in == 338) begin
					state<=2;
					out<=120;
				end
				if(in == 339) begin
					state<=2;
					out<=121;
				end
				if(in == 340) begin
					state<=2;
					out<=122;
				end
				if(in == 341) begin
					state<=2;
					out<=123;
				end
				if(in == 342) begin
					state<=2;
					out<=124;
				end
				if(in == 343) begin
					state<=2;
					out<=125;
				end
				if(in == 344) begin
					state<=2;
					out<=126;
				end
				if(in == 345) begin
					state<=2;
					out<=127;
				end
				if(in == 346) begin
					state<=2;
					out<=128;
				end
				if(in == 347) begin
					state<=2;
					out<=129;
				end
				if(in == 348) begin
					state<=2;
					out<=130;
				end
				if(in == 349) begin
					state<=3;
					out<=131;
				end
				if(in == 350) begin
					state<=6;
					out<=132;
				end
				if(in == 351) begin
					state<=3;
					out<=133;
				end
				if(in == 352) begin
					state<=7;
					out<=134;
				end
				if(in == 353) begin
					state<=3;
					out<=135;
				end
				if(in == 354) begin
					state<=7;
					out<=136;
				end
				if(in == 355) begin
					state<=7;
					out<=137;
				end
				if(in == 356) begin
					state<=7;
					out<=138;
				end
				if(in == 357) begin
					state<=7;
					out<=139;
				end
				if(in == 358) begin
					state<=7;
					out<=140;
				end
				if(in == 359) begin
					state<=7;
					out<=141;
				end
				if(in == 360) begin
					state<=7;
					out<=142;
				end
				if(in == 361) begin
					state<=7;
					out<=143;
				end
				if(in == 362) begin
					state<=7;
					out<=144;
				end
				if(in == 363) begin
					state<=7;
					out<=145;
				end
				if(in == 364) begin
					state<=7;
					out<=146;
				end
				if(in == 365) begin
					state<=7;
					out<=147;
				end
				if(in == 366) begin
					state<=7;
					out<=148;
				end
				if(in == 367) begin
					state<=7;
					out<=149;
				end
				if(in == 368) begin
					state<=7;
					out<=150;
				end
				if(in == 369) begin
					state<=7;
					out<=151;
				end
				if(in == 370) begin
					state<=7;
					out<=152;
				end
				if(in == 371) begin
					state<=7;
					out<=153;
				end
				if(in == 372) begin
					state<=7;
					out<=154;
				end
				if(in == 373) begin
					state<=7;
					out<=155;
				end
				if(in == 374) begin
					state<=7;
					out<=156;
				end
				if(in == 375) begin
					state<=7;
					out<=157;
				end
				if(in == 376) begin
					state<=7;
					out<=158;
				end
				if(in == 377) begin
					state<=7;
					out<=159;
				end
				if(in == 378) begin
					state<=7;
					out<=160;
				end
				if(in == 379) begin
					state<=7;
					out<=161;
				end
				if(in == 380) begin
					state<=7;
					out<=162;
				end
				if(in == 381) begin
					state<=7;
					out<=163;
				end
				if(in == 382) begin
					state<=7;
					out<=164;
				end
				if(in == 383) begin
					state<=7;
					out<=165;
				end
				if(in == 384) begin
					state<=7;
					out<=166;
				end
				if(in == 385) begin
					state<=7;
					out<=167;
				end
				if(in == 386) begin
					state<=7;
					out<=168;
				end
				if(in == 387) begin
					state<=7;
					out<=169;
				end
				if(in == 388) begin
					state<=7;
					out<=170;
				end
				if(in == 389) begin
					state<=7;
					out<=171;
				end
				if(in == 390) begin
					state<=7;
					out<=172;
				end
				if(in == 391) begin
					state<=7;
					out<=173;
				end
				if(in == 392) begin
					state<=7;
					out<=174;
				end
				if(in == 393) begin
					state<=7;
					out<=175;
				end
				if(in == 394) begin
					state<=7;
					out<=176;
				end
				if(in == 395) begin
					state<=7;
					out<=177;
				end
				if(in == 396) begin
					state<=7;
					out<=178;
				end
				if(in == 397) begin
					state<=7;
					out<=179;
				end
				if(in == 398) begin
					state<=7;
					out<=180;
				end
				if(in == 399) begin
					state<=7;
					out<=181;
				end
				if(in == 400) begin
					state<=7;
					out<=182;
				end
				if(in == 401) begin
					state<=3;
					out<=183;
				end
				if(in == 402) begin
					state<=6;
					out<=184;
				end
				if(in == 403) begin
					state<=3;
					out<=185;
				end
				if(in == 404) begin
					state<=7;
					out<=186;
				end
				if(in == 405) begin
					state<=3;
					out<=187;
				end
				if(in == 406) begin
					state<=7;
					out<=188;
				end
				if(in == 407) begin
					state<=7;
					out<=189;
				end
				if(in == 408) begin
					state<=7;
					out<=190;
				end
				if(in == 409) begin
					state<=7;
					out<=191;
				end
				if(in == 410) begin
					state<=7;
					out<=192;
				end
				if(in == 411) begin
					state<=7;
					out<=193;
				end
				if(in == 412) begin
					state<=7;
					out<=194;
				end
				if(in == 413) begin
					state<=7;
					out<=195;
				end
				if(in == 414) begin
					state<=7;
					out<=196;
				end
				if(in == 415) begin
					state<=7;
					out<=197;
				end
				if(in == 416) begin
					state<=7;
					out<=198;
				end
				if(in == 417) begin
					state<=7;
					out<=199;
				end
				if(in == 418) begin
					state<=7;
					out<=200;
				end
				if(in == 419) begin
					state<=7;
					out<=201;
				end
				if(in == 420) begin
					state<=7;
					out<=202;
				end
				if(in == 421) begin
					state<=7;
					out<=203;
				end
				if(in == 422) begin
					state<=7;
					out<=204;
				end
				if(in == 423) begin
					state<=7;
					out<=205;
				end
				if(in == 424) begin
					state<=7;
					out<=206;
				end
				if(in == 425) begin
					state<=7;
					out<=207;
				end
				if(in == 426) begin
					state<=7;
					out<=208;
				end
				if(in == 427) begin
					state<=7;
					out<=209;
				end
				if(in == 428) begin
					state<=7;
					out<=210;
				end
				if(in == 429) begin
					state<=7;
					out<=211;
				end
				if(in == 430) begin
					state<=7;
					out<=212;
				end
				if(in == 431) begin
					state<=7;
					out<=213;
				end
				if(in == 432) begin
					state<=7;
					out<=214;
				end
				if(in == 433) begin
					state<=7;
					out<=215;
				end
				if(in == 434) begin
					state<=7;
					out<=216;
				end
				if(in == 435) begin
					state<=7;
					out<=217;
				end
				if(in == 436) begin
					state<=7;
					out<=218;
				end
				if(in == 437) begin
					state<=7;
					out<=219;
				end
				if(in == 438) begin
					state<=7;
					out<=220;
				end
				if(in == 439) begin
					state<=7;
					out<=221;
				end
				if(in == 440) begin
					state<=7;
					out<=222;
				end
				if(in == 441) begin
					state<=7;
					out<=223;
				end
				if(in == 442) begin
					state<=7;
					out<=224;
				end
				if(in == 443) begin
					state<=7;
					out<=225;
				end
				if(in == 444) begin
					state<=7;
					out<=226;
				end
				if(in == 445) begin
					state<=7;
					out<=227;
				end
				if(in == 446) begin
					state<=7;
					out<=228;
				end
				if(in == 447) begin
					state<=7;
					out<=229;
				end
				if(in == 448) begin
					state<=7;
					out<=230;
				end
				if(in == 449) begin
					state<=7;
					out<=231;
				end
				if(in == 450) begin
					state<=7;
					out<=232;
				end
				if(in == 451) begin
					state<=7;
					out<=233;
				end
				if(in == 452) begin
					state<=7;
					out<=234;
				end
				if(in == 453) begin
					state<=2;
					out<=235;
				end
				if(in == 454) begin
					state<=2;
					out<=236;
				end
				if(in == 455) begin
					state<=2;
					out<=237;
				end
				if(in == 456) begin
					state<=2;
					out<=238;
				end
				if(in == 457) begin
					state<=2;
					out<=239;
				end
				if(in == 458) begin
					state<=2;
					out<=240;
				end
				if(in == 459) begin
					state<=2;
					out<=241;
				end
				if(in == 460) begin
					state<=2;
					out<=242;
				end
				if(in == 461) begin
					state<=2;
					out<=243;
				end
				if(in == 462) begin
					state<=2;
					out<=244;
				end
				if(in == 463) begin
					state<=2;
					out<=245;
				end
				if(in == 464) begin
					state<=2;
					out<=246;
				end
				if(in == 465) begin
					state<=3;
					out<=247;
				end
				if(in == 466) begin
					state<=6;
					out<=248;
				end
				if(in == 467) begin
					state<=3;
					out<=249;
				end
				if(in == 468) begin
					state<=7;
					out<=250;
				end
				if(in == 469) begin
					state<=3;
					out<=251;
				end
				if(in == 470) begin
					state<=7;
					out<=252;
				end
				if(in == 471) begin
					state<=7;
					out<=253;
				end
				if(in == 472) begin
					state<=7;
					out<=254;
				end
				if(in == 473) begin
					state<=7;
					out<=255;
				end
				if(in == 474) begin
					state<=7;
					out<=0;
				end
				if(in == 475) begin
					state<=7;
					out<=1;
				end
				if(in == 476) begin
					state<=7;
					out<=2;
				end
				if(in == 477) begin
					state<=7;
					out<=3;
				end
				if(in == 478) begin
					state<=7;
					out<=4;
				end
				if(in == 479) begin
					state<=7;
					out<=5;
				end
				if(in == 480) begin
					state<=7;
					out<=6;
				end
				if(in == 481) begin
					state<=7;
					out<=7;
				end
				if(in == 482) begin
					state<=7;
					out<=8;
				end
				if(in == 483) begin
					state<=7;
					out<=9;
				end
				if(in == 484) begin
					state<=7;
					out<=10;
				end
				if(in == 485) begin
					state<=7;
					out<=11;
				end
				if(in == 486) begin
					state<=7;
					out<=12;
				end
				if(in == 487) begin
					state<=7;
					out<=13;
				end
				if(in == 488) begin
					state<=7;
					out<=14;
				end
				if(in == 489) begin
					state<=7;
					out<=15;
				end
				if(in == 490) begin
					state<=7;
					out<=16;
				end
				if(in == 491) begin
					state<=7;
					out<=17;
				end
				if(in == 492) begin
					state<=7;
					out<=18;
				end
				if(in == 493) begin
					state<=7;
					out<=19;
				end
				if(in == 494) begin
					state<=7;
					out<=20;
				end
				if(in == 495) begin
					state<=7;
					out<=21;
				end
				if(in == 496) begin
					state<=7;
					out<=22;
				end
				if(in == 497) begin
					state<=7;
					out<=23;
				end
				if(in == 498) begin
					state<=7;
					out<=24;
				end
				if(in == 499) begin
					state<=7;
					out<=25;
				end
				if(in == 500) begin
					state<=7;
					out<=26;
				end
				if(in == 501) begin
					state<=7;
					out<=27;
				end
				if(in == 502) begin
					state<=7;
					out<=28;
				end
				if(in == 503) begin
					state<=7;
					out<=29;
				end
				if(in == 504) begin
					state<=7;
					out<=30;
				end
				if(in == 505) begin
					state<=7;
					out<=31;
				end
				if(in == 506) begin
					state<=7;
					out<=32;
				end
				if(in == 507) begin
					state<=7;
					out<=33;
				end
				if(in == 508) begin
					state<=7;
					out<=34;
				end
				if(in == 509) begin
					state<=7;
					out<=35;
				end
				if(in == 510) begin
					state<=7;
					out<=36;
				end
				if(in == 511) begin
					state<=7;
					out<=37;
				end
				if(in == 512) begin
					state<=7;
					out<=38;
				end
				if(in == 513) begin
					state<=7;
					out<=39;
				end
				if(in == 514) begin
					state<=7;
					out<=40;
				end
				if(in == 515) begin
					state<=7;
					out<=41;
				end
				if(in == 516) begin
					state<=7;
					out<=42;
				end
				if(in == 517) begin
					state<=3;
					out<=43;
				end
				if(in == 518) begin
					state<=6;
					out<=44;
				end
				if(in == 519) begin
					state<=3;
					out<=45;
				end
				if(in == 520) begin
					state<=7;
					out<=46;
				end
				if(in == 521) begin
					state<=3;
					out<=47;
				end
				if(in == 522) begin
					state<=7;
					out<=48;
				end
				if(in == 523) begin
					state<=7;
					out<=49;
				end
				if(in == 524) begin
					state<=7;
					out<=50;
				end
				if(in == 525) begin
					state<=7;
					out<=51;
				end
				if(in == 526) begin
					state<=7;
					out<=52;
				end
				if(in == 527) begin
					state<=7;
					out<=53;
				end
				if(in == 528) begin
					state<=7;
					out<=54;
				end
				if(in == 529) begin
					state<=7;
					out<=55;
				end
				if(in == 530) begin
					state<=7;
					out<=56;
				end
				if(in == 531) begin
					state<=7;
					out<=57;
				end
				if(in == 532) begin
					state<=7;
					out<=58;
				end
				if(in == 533) begin
					state<=7;
					out<=59;
				end
				if(in == 534) begin
					state<=7;
					out<=60;
				end
				if(in == 535) begin
					state<=7;
					out<=61;
				end
				if(in == 536) begin
					state<=7;
					out<=62;
				end
				if(in == 537) begin
					state<=7;
					out<=63;
				end
				if(in == 538) begin
					state<=7;
					out<=64;
				end
				if(in == 539) begin
					state<=7;
					out<=65;
				end
				if(in == 540) begin
					state<=7;
					out<=66;
				end
				if(in == 541) begin
					state<=7;
					out<=67;
				end
				if(in == 542) begin
					state<=7;
					out<=68;
				end
				if(in == 543) begin
					state<=7;
					out<=69;
				end
				if(in == 544) begin
					state<=7;
					out<=70;
				end
				if(in == 545) begin
					state<=7;
					out<=71;
				end
				if(in == 546) begin
					state<=7;
					out<=72;
				end
				if(in == 547) begin
					state<=7;
					out<=73;
				end
				if(in == 548) begin
					state<=7;
					out<=74;
				end
				if(in == 549) begin
					state<=7;
					out<=75;
				end
				if(in == 550) begin
					state<=7;
					out<=76;
				end
				if(in == 551) begin
					state<=7;
					out<=77;
				end
				if(in == 552) begin
					state<=7;
					out<=78;
				end
				if(in == 553) begin
					state<=7;
					out<=79;
				end
				if(in == 554) begin
					state<=7;
					out<=80;
				end
				if(in == 555) begin
					state<=7;
					out<=81;
				end
				if(in == 556) begin
					state<=7;
					out<=82;
				end
				if(in == 557) begin
					state<=7;
					out<=83;
				end
				if(in == 558) begin
					state<=7;
					out<=84;
				end
				if(in == 559) begin
					state<=7;
					out<=85;
				end
				if(in == 560) begin
					state<=7;
					out<=86;
				end
				if(in == 561) begin
					state<=7;
					out<=87;
				end
				if(in == 562) begin
					state<=7;
					out<=88;
				end
				if(in == 563) begin
					state<=7;
					out<=89;
				end
				if(in == 564) begin
					state<=7;
					out<=90;
				end
				if(in == 565) begin
					state<=7;
					out<=91;
				end
				if(in == 566) begin
					state<=7;
					out<=92;
				end
				if(in == 567) begin
					state<=7;
					out<=93;
				end
				if(in == 568) begin
					state<=7;
					out<=94;
				end
				if(in == 569) begin
					state<=2;
					out<=95;
				end
				if(in == 570) begin
					state<=2;
					out<=96;
				end
				if(in == 571) begin
					state<=2;
					out<=97;
				end
				if(in == 572) begin
					state<=2;
					out<=98;
				end
				if(in == 573) begin
					state<=2;
					out<=99;
				end
				if(in == 574) begin
					state<=2;
					out<=100;
				end
				if(in == 575) begin
					state<=2;
					out<=101;
				end
				if(in == 576) begin
					state<=2;
					out<=102;
				end
				if(in == 577) begin
					state<=2;
					out<=103;
				end
				if(in == 578) begin
					state<=2;
					out<=104;
				end
				if(in == 579) begin
					state<=2;
					out<=105;
				end
				if(in == 580) begin
					state<=2;
					out<=106;
				end
				if(in == 581) begin
					state<=3;
					out<=107;
				end
				if(in == 582) begin
					state<=6;
					out<=108;
				end
				if(in == 583) begin
					state<=3;
					out<=109;
				end
				if(in == 584) begin
					state<=7;
					out<=110;
				end
				if(in == 585) begin
					state<=3;
					out<=111;
				end
				if(in == 586) begin
					state<=7;
					out<=112;
				end
				if(in == 587) begin
					state<=7;
					out<=113;
				end
				if(in == 588) begin
					state<=7;
					out<=114;
				end
				if(in == 589) begin
					state<=7;
					out<=115;
				end
				if(in == 590) begin
					state<=7;
					out<=116;
				end
				if(in == 591) begin
					state<=7;
					out<=117;
				end
				if(in == 592) begin
					state<=7;
					out<=118;
				end
				if(in == 593) begin
					state<=7;
					out<=119;
				end
				if(in == 594) begin
					state<=7;
					out<=120;
				end
				if(in == 595) begin
					state<=7;
					out<=121;
				end
				if(in == 596) begin
					state<=7;
					out<=122;
				end
				if(in == 597) begin
					state<=7;
					out<=123;
				end
				if(in == 598) begin
					state<=7;
					out<=124;
				end
				if(in == 599) begin
					state<=7;
					out<=125;
				end
				if(in == 600) begin
					state<=7;
					out<=126;
				end
				if(in == 601) begin
					state<=7;
					out<=127;
				end
				if(in == 602) begin
					state<=7;
					out<=128;
				end
				if(in == 603) begin
					state<=7;
					out<=129;
				end
				if(in == 604) begin
					state<=7;
					out<=130;
				end
				if(in == 605) begin
					state<=7;
					out<=131;
				end
				if(in == 606) begin
					state<=7;
					out<=132;
				end
				if(in == 607) begin
					state<=7;
					out<=133;
				end
				if(in == 608) begin
					state<=7;
					out<=134;
				end
				if(in == 609) begin
					state<=7;
					out<=135;
				end
				if(in == 610) begin
					state<=7;
					out<=136;
				end
				if(in == 611) begin
					state<=7;
					out<=137;
				end
				if(in == 612) begin
					state<=7;
					out<=138;
				end
				if(in == 613) begin
					state<=7;
					out<=139;
				end
				if(in == 614) begin
					state<=7;
					out<=140;
				end
				if(in == 615) begin
					state<=7;
					out<=141;
				end
				if(in == 616) begin
					state<=7;
					out<=142;
				end
				if(in == 617) begin
					state<=7;
					out<=143;
				end
				if(in == 618) begin
					state<=7;
					out<=144;
				end
				if(in == 619) begin
					state<=7;
					out<=145;
				end
				if(in == 620) begin
					state<=7;
					out<=146;
				end
				if(in == 621) begin
					state<=7;
					out<=147;
				end
				if(in == 622) begin
					state<=7;
					out<=148;
				end
				if(in == 623) begin
					state<=7;
					out<=149;
				end
				if(in == 624) begin
					state<=7;
					out<=150;
				end
				if(in == 625) begin
					state<=7;
					out<=151;
				end
				if(in == 626) begin
					state<=7;
					out<=152;
				end
				if(in == 627) begin
					state<=7;
					out<=153;
				end
				if(in == 628) begin
					state<=7;
					out<=154;
				end
				if(in == 629) begin
					state<=7;
					out<=155;
				end
				if(in == 630) begin
					state<=7;
					out<=156;
				end
				if(in == 631) begin
					state<=7;
					out<=157;
				end
				if(in == 632) begin
					state<=7;
					out<=158;
				end
				if(in == 633) begin
					state<=3;
					out<=159;
				end
				if(in == 634) begin
					state<=6;
					out<=160;
				end
				if(in == 635) begin
					state<=3;
					out<=161;
				end
				if(in == 636) begin
					state<=7;
					out<=162;
				end
				if(in == 637) begin
					state<=3;
					out<=163;
				end
				if(in == 638) begin
					state<=7;
					out<=164;
				end
				if(in == 639) begin
					state<=7;
					out<=165;
				end
				if(in == 640) begin
					state<=7;
					out<=166;
				end
				if(in == 641) begin
					state<=7;
					out<=167;
				end
				if(in == 642) begin
					state<=7;
					out<=168;
				end
				if(in == 643) begin
					state<=7;
					out<=169;
				end
				if(in == 644) begin
					state<=7;
					out<=170;
				end
				if(in == 645) begin
					state<=7;
					out<=171;
				end
				if(in == 646) begin
					state<=7;
					out<=172;
				end
				if(in == 647) begin
					state<=7;
					out<=173;
				end
				if(in == 648) begin
					state<=7;
					out<=174;
				end
				if(in == 649) begin
					state<=7;
					out<=175;
				end
				if(in == 650) begin
					state<=7;
					out<=176;
				end
				if(in == 651) begin
					state<=7;
					out<=177;
				end
				if(in == 652) begin
					state<=7;
					out<=178;
				end
				if(in == 653) begin
					state<=7;
					out<=179;
				end
				if(in == 654) begin
					state<=7;
					out<=180;
				end
				if(in == 655) begin
					state<=7;
					out<=181;
				end
				if(in == 656) begin
					state<=7;
					out<=182;
				end
				if(in == 657) begin
					state<=7;
					out<=183;
				end
				if(in == 658) begin
					state<=7;
					out<=184;
				end
				if(in == 659) begin
					state<=7;
					out<=185;
				end
				if(in == 660) begin
					state<=7;
					out<=186;
				end
				if(in == 661) begin
					state<=7;
					out<=187;
				end
				if(in == 662) begin
					state<=7;
					out<=188;
				end
				if(in == 663) begin
					state<=7;
					out<=189;
				end
				if(in == 664) begin
					state<=7;
					out<=190;
				end
				if(in == 665) begin
					state<=7;
					out<=191;
				end
				if(in == 666) begin
					state<=7;
					out<=192;
				end
				if(in == 667) begin
					state<=7;
					out<=193;
				end
				if(in == 668) begin
					state<=7;
					out<=194;
				end
				if(in == 669) begin
					state<=7;
					out<=195;
				end
				if(in == 670) begin
					state<=7;
					out<=196;
				end
				if(in == 671) begin
					state<=7;
					out<=197;
				end
				if(in == 672) begin
					state<=7;
					out<=198;
				end
				if(in == 673) begin
					state<=7;
					out<=199;
				end
				if(in == 674) begin
					state<=7;
					out<=200;
				end
				if(in == 675) begin
					state<=7;
					out<=201;
				end
				if(in == 676) begin
					state<=7;
					out<=202;
				end
				if(in == 677) begin
					state<=7;
					out<=203;
				end
				if(in == 678) begin
					state<=7;
					out<=204;
				end
				if(in == 679) begin
					state<=7;
					out<=205;
				end
				if(in == 680) begin
					state<=7;
					out<=206;
				end
				if(in == 681) begin
					state<=7;
					out<=207;
				end
				if(in == 682) begin
					state<=7;
					out<=208;
				end
				if(in == 683) begin
					state<=7;
					out<=209;
				end
				if(in == 684) begin
					state<=7;
					out<=210;
				end
				if(in == 685) begin
					state<=2;
					out<=211;
				end
				if(in == 686) begin
					state<=2;
					out<=212;
				end
				if(in == 687) begin
					state<=2;
					out<=213;
				end
				if(in == 688) begin
					state<=2;
					out<=214;
				end
				if(in == 689) begin
					state<=2;
					out<=215;
				end
				if(in == 690) begin
					state<=2;
					out<=216;
				end
				if(in == 691) begin
					state<=2;
					out<=217;
				end
				if(in == 692) begin
					state<=2;
					out<=218;
				end
				if(in == 693) begin
					state<=2;
					out<=219;
				end
				if(in == 694) begin
					state<=2;
					out<=220;
				end
				if(in == 695) begin
					state<=2;
					out<=221;
				end
				if(in == 696) begin
					state<=2;
					out<=222;
				end
				if(in == 697) begin
					state<=3;
					out<=223;
				end
				if(in == 698) begin
					state<=6;
					out<=224;
				end
				if(in == 699) begin
					state<=3;
					out<=225;
				end
				if(in == 700) begin
					state<=7;
					out<=226;
				end
				if(in == 701) begin
					state<=3;
					out<=227;
				end
				if(in == 702) begin
					state<=7;
					out<=228;
				end
				if(in == 703) begin
					state<=7;
					out<=229;
				end
				if(in == 704) begin
					state<=7;
					out<=230;
				end
				if(in == 705) begin
					state<=7;
					out<=231;
				end
				if(in == 706) begin
					state<=7;
					out<=232;
				end
				if(in == 707) begin
					state<=7;
					out<=233;
				end
				if(in == 708) begin
					state<=7;
					out<=234;
				end
				if(in == 709) begin
					state<=7;
					out<=235;
				end
				if(in == 710) begin
					state<=7;
					out<=236;
				end
				if(in == 711) begin
					state<=7;
					out<=237;
				end
				if(in == 712) begin
					state<=7;
					out<=238;
				end
				if(in == 713) begin
					state<=7;
					out<=239;
				end
				if(in == 714) begin
					state<=7;
					out<=240;
				end
				if(in == 715) begin
					state<=7;
					out<=241;
				end
				if(in == 716) begin
					state<=7;
					out<=242;
				end
				if(in == 717) begin
					state<=7;
					out<=243;
				end
				if(in == 718) begin
					state<=7;
					out<=244;
				end
				if(in == 719) begin
					state<=7;
					out<=245;
				end
				if(in == 720) begin
					state<=7;
					out<=246;
				end
				if(in == 721) begin
					state<=7;
					out<=247;
				end
				if(in == 722) begin
					state<=7;
					out<=248;
				end
				if(in == 723) begin
					state<=7;
					out<=249;
				end
				if(in == 724) begin
					state<=7;
					out<=250;
				end
				if(in == 725) begin
					state<=7;
					out<=251;
				end
				if(in == 726) begin
					state<=7;
					out<=252;
				end
				if(in == 727) begin
					state<=7;
					out<=253;
				end
				if(in == 728) begin
					state<=7;
					out<=254;
				end
				if(in == 729) begin
					state<=7;
					out<=255;
				end
				if(in == 730) begin
					state<=7;
					out<=0;
				end
				if(in == 731) begin
					state<=7;
					out<=1;
				end
				if(in == 732) begin
					state<=7;
					out<=2;
				end
				if(in == 733) begin
					state<=7;
					out<=3;
				end
				if(in == 734) begin
					state<=7;
					out<=4;
				end
				if(in == 735) begin
					state<=7;
					out<=5;
				end
				if(in == 736) begin
					state<=7;
					out<=6;
				end
				if(in == 737) begin
					state<=7;
					out<=7;
				end
				if(in == 738) begin
					state<=7;
					out<=8;
				end
				if(in == 739) begin
					state<=7;
					out<=9;
				end
				if(in == 740) begin
					state<=7;
					out<=10;
				end
				if(in == 741) begin
					state<=7;
					out<=11;
				end
				if(in == 742) begin
					state<=7;
					out<=12;
				end
				if(in == 743) begin
					state<=7;
					out<=13;
				end
				if(in == 744) begin
					state<=7;
					out<=14;
				end
				if(in == 745) begin
					state<=7;
					out<=15;
				end
				if(in == 746) begin
					state<=7;
					out<=16;
				end
				if(in == 747) begin
					state<=7;
					out<=17;
				end
				if(in == 748) begin
					state<=7;
					out<=18;
				end
				if(in == 749) begin
					state<=3;
					out<=19;
				end
				if(in == 750) begin
					state<=6;
					out<=20;
				end
				if(in == 751) begin
					state<=3;
					out<=21;
				end
				if(in == 752) begin
					state<=7;
					out<=22;
				end
				if(in == 753) begin
					state<=3;
					out<=23;
				end
				if(in == 754) begin
					state<=7;
					out<=24;
				end
				if(in == 755) begin
					state<=7;
					out<=25;
				end
				if(in == 756) begin
					state<=7;
					out<=26;
				end
				if(in == 757) begin
					state<=7;
					out<=27;
				end
				if(in == 758) begin
					state<=7;
					out<=28;
				end
				if(in == 759) begin
					state<=7;
					out<=29;
				end
				if(in == 760) begin
					state<=7;
					out<=30;
				end
				if(in == 761) begin
					state<=7;
					out<=31;
				end
				if(in == 762) begin
					state<=7;
					out<=32;
				end
				if(in == 763) begin
					state<=7;
					out<=33;
				end
				if(in == 764) begin
					state<=7;
					out<=34;
				end
				if(in == 765) begin
					state<=7;
					out<=35;
				end
				if(in == 766) begin
					state<=7;
					out<=36;
				end
				if(in == 767) begin
					state<=7;
					out<=37;
				end
				if(in == 768) begin
					state<=7;
					out<=38;
				end
				if(in == 769) begin
					state<=7;
					out<=39;
				end
				if(in == 770) begin
					state<=7;
					out<=40;
				end
				if(in == 771) begin
					state<=7;
					out<=41;
				end
				if(in == 772) begin
					state<=7;
					out<=42;
				end
				if(in == 773) begin
					state<=7;
					out<=43;
				end
				if(in == 774) begin
					state<=7;
					out<=44;
				end
				if(in == 775) begin
					state<=7;
					out<=45;
				end
				if(in == 776) begin
					state<=7;
					out<=46;
				end
				if(in == 777) begin
					state<=7;
					out<=47;
				end
				if(in == 778) begin
					state<=7;
					out<=48;
				end
				if(in == 779) begin
					state<=7;
					out<=49;
				end
				if(in == 780) begin
					state<=7;
					out<=50;
				end
				if(in == 781) begin
					state<=7;
					out<=51;
				end
				if(in == 782) begin
					state<=7;
					out<=52;
				end
				if(in == 783) begin
					state<=7;
					out<=53;
				end
				if(in == 784) begin
					state<=7;
					out<=54;
				end
				if(in == 785) begin
					state<=7;
					out<=55;
				end
				if(in == 786) begin
					state<=7;
					out<=56;
				end
				if(in == 787) begin
					state<=7;
					out<=57;
				end
				if(in == 788) begin
					state<=7;
					out<=58;
				end
				if(in == 789) begin
					state<=7;
					out<=59;
				end
				if(in == 790) begin
					state<=7;
					out<=60;
				end
				if(in == 791) begin
					state<=7;
					out<=61;
				end
				if(in == 792) begin
					state<=7;
					out<=62;
				end
				if(in == 793) begin
					state<=7;
					out<=63;
				end
				if(in == 794) begin
					state<=7;
					out<=64;
				end
				if(in == 795) begin
					state<=7;
					out<=65;
				end
				if(in == 796) begin
					state<=7;
					out<=66;
				end
				if(in == 797) begin
					state<=7;
					out<=67;
				end
				if(in == 798) begin
					state<=7;
					out<=68;
				end
				if(in == 799) begin
					state<=7;
					out<=69;
				end
				if(in == 800) begin
					state<=7;
					out<=70;
				end
				if(in == 801) begin
					state<=2;
					out<=71;
				end
				if(in == 802) begin
					state<=2;
					out<=72;
				end
				if(in == 803) begin
					state<=2;
					out<=73;
				end
				if(in == 804) begin
					state<=2;
					out<=74;
				end
				if(in == 805) begin
					state<=2;
					out<=75;
				end
				if(in == 806) begin
					state<=2;
					out<=76;
				end
				if(in == 807) begin
					state<=2;
					out<=77;
				end
				if(in == 808) begin
					state<=2;
					out<=78;
				end
				if(in == 809) begin
					state<=2;
					out<=79;
				end
				if(in == 810) begin
					state<=2;
					out<=80;
				end
				if(in == 811) begin
					state<=2;
					out<=81;
				end
				if(in == 812) begin
					state<=2;
					out<=82;
				end
				if(in == 813) begin
					state<=3;
					out<=83;
				end
				if(in == 814) begin
					state<=6;
					out<=84;
				end
				if(in == 815) begin
					state<=3;
					out<=85;
				end
				if(in == 816) begin
					state<=7;
					out<=86;
				end
				if(in == 817) begin
					state<=3;
					out<=87;
				end
				if(in == 818) begin
					state<=7;
					out<=88;
				end
				if(in == 819) begin
					state<=7;
					out<=89;
				end
				if(in == 820) begin
					state<=7;
					out<=90;
				end
				if(in == 821) begin
					state<=7;
					out<=91;
				end
				if(in == 822) begin
					state<=7;
					out<=92;
				end
				if(in == 823) begin
					state<=7;
					out<=93;
				end
				if(in == 824) begin
					state<=7;
					out<=94;
				end
				if(in == 825) begin
					state<=7;
					out<=95;
				end
				if(in == 826) begin
					state<=7;
					out<=96;
				end
				if(in == 827) begin
					state<=7;
					out<=97;
				end
				if(in == 828) begin
					state<=7;
					out<=98;
				end
				if(in == 829) begin
					state<=7;
					out<=99;
				end
				if(in == 830) begin
					state<=7;
					out<=100;
				end
				if(in == 831) begin
					state<=7;
					out<=101;
				end
				if(in == 832) begin
					state<=7;
					out<=102;
				end
				if(in == 833) begin
					state<=7;
					out<=103;
				end
				if(in == 834) begin
					state<=7;
					out<=104;
				end
				if(in == 835) begin
					state<=7;
					out<=105;
				end
				if(in == 836) begin
					state<=7;
					out<=106;
				end
				if(in == 837) begin
					state<=7;
					out<=107;
				end
				if(in == 838) begin
					state<=7;
					out<=108;
				end
				if(in == 839) begin
					state<=7;
					out<=109;
				end
				if(in == 840) begin
					state<=7;
					out<=110;
				end
				if(in == 841) begin
					state<=7;
					out<=111;
				end
				if(in == 842) begin
					state<=7;
					out<=112;
				end
				if(in == 843) begin
					state<=7;
					out<=113;
				end
				if(in == 844) begin
					state<=7;
					out<=114;
				end
				if(in == 845) begin
					state<=7;
					out<=115;
				end
				if(in == 846) begin
					state<=7;
					out<=116;
				end
				if(in == 847) begin
					state<=7;
					out<=117;
				end
				if(in == 848) begin
					state<=7;
					out<=118;
				end
				if(in == 849) begin
					state<=7;
					out<=119;
				end
				if(in == 850) begin
					state<=7;
					out<=120;
				end
				if(in == 851) begin
					state<=7;
					out<=121;
				end
				if(in == 852) begin
					state<=7;
					out<=122;
				end
				if(in == 853) begin
					state<=7;
					out<=123;
				end
				if(in == 854) begin
					state<=7;
					out<=124;
				end
				if(in == 855) begin
					state<=7;
					out<=125;
				end
				if(in == 856) begin
					state<=7;
					out<=126;
				end
				if(in == 857) begin
					state<=7;
					out<=127;
				end
				if(in == 858) begin
					state<=7;
					out<=128;
				end
				if(in == 859) begin
					state<=7;
					out<=129;
				end
				if(in == 860) begin
					state<=7;
					out<=130;
				end
				if(in == 861) begin
					state<=7;
					out<=131;
				end
				if(in == 862) begin
					state<=7;
					out<=132;
				end
				if(in == 863) begin
					state<=7;
					out<=133;
				end
				if(in == 864) begin
					state<=7;
					out<=134;
				end
				if(in == 865) begin
					state<=3;
					out<=135;
				end
				if(in == 866) begin
					state<=6;
					out<=136;
				end
				if(in == 867) begin
					state<=3;
					out<=137;
				end
				if(in == 868) begin
					state<=7;
					out<=138;
				end
				if(in == 869) begin
					state<=3;
					out<=139;
				end
				if(in == 870) begin
					state<=7;
					out<=140;
				end
				if(in == 871) begin
					state<=7;
					out<=141;
				end
				if(in == 872) begin
					state<=7;
					out<=142;
				end
				if(in == 873) begin
					state<=7;
					out<=143;
				end
				if(in == 874) begin
					state<=7;
					out<=144;
				end
				if(in == 875) begin
					state<=7;
					out<=145;
				end
				if(in == 876) begin
					state<=7;
					out<=146;
				end
				if(in == 877) begin
					state<=7;
					out<=147;
				end
				if(in == 878) begin
					state<=7;
					out<=148;
				end
				if(in == 879) begin
					state<=7;
					out<=149;
				end
				if(in == 880) begin
					state<=7;
					out<=150;
				end
				if(in == 881) begin
					state<=7;
					out<=151;
				end
				if(in == 882) begin
					state<=7;
					out<=152;
				end
				if(in == 883) begin
					state<=7;
					out<=153;
				end
				if(in == 884) begin
					state<=7;
					out<=154;
				end
				if(in == 885) begin
					state<=7;
					out<=155;
				end
				if(in == 886) begin
					state<=7;
					out<=156;
				end
				if(in == 887) begin
					state<=7;
					out<=157;
				end
				if(in == 888) begin
					state<=7;
					out<=158;
				end
				if(in == 889) begin
					state<=7;
					out<=159;
				end
				if(in == 890) begin
					state<=7;
					out<=160;
				end
				if(in == 891) begin
					state<=7;
					out<=161;
				end
				if(in == 892) begin
					state<=7;
					out<=162;
				end
				if(in == 893) begin
					state<=7;
					out<=163;
				end
				if(in == 894) begin
					state<=7;
					out<=164;
				end
				if(in == 895) begin
					state<=7;
					out<=165;
				end
				if(in == 896) begin
					state<=7;
					out<=166;
				end
				if(in == 897) begin
					state<=7;
					out<=167;
				end
				if(in == 898) begin
					state<=7;
					out<=168;
				end
				if(in == 899) begin
					state<=7;
					out<=169;
				end
				if(in == 900) begin
					state<=7;
					out<=170;
				end
				if(in == 901) begin
					state<=7;
					out<=171;
				end
				if(in == 902) begin
					state<=7;
					out<=172;
				end
				if(in == 903) begin
					state<=7;
					out<=173;
				end
				if(in == 904) begin
					state<=7;
					out<=174;
				end
				if(in == 905) begin
					state<=7;
					out<=175;
				end
				if(in == 906) begin
					state<=7;
					out<=176;
				end
				if(in == 907) begin
					state<=7;
					out<=177;
				end
				if(in == 908) begin
					state<=7;
					out<=178;
				end
				if(in == 909) begin
					state<=7;
					out<=179;
				end
				if(in == 910) begin
					state<=7;
					out<=180;
				end
				if(in == 911) begin
					state<=7;
					out<=181;
				end
				if(in == 912) begin
					state<=7;
					out<=182;
				end
				if(in == 913) begin
					state<=7;
					out<=183;
				end
				if(in == 914) begin
					state<=7;
					out<=184;
				end
				if(in == 915) begin
					state<=7;
					out<=185;
				end
				if(in == 916) begin
					state<=7;
					out<=186;
				end
				if(in == 917) begin
					state<=2;
					out<=187;
				end
				if(in == 918) begin
					state<=2;
					out<=188;
				end
				if(in == 919) begin
					state<=2;
					out<=189;
				end
				if(in == 920) begin
					state<=2;
					out<=190;
				end
				if(in == 921) begin
					state<=2;
					out<=191;
				end
				if(in == 922) begin
					state<=2;
					out<=192;
				end
				if(in == 923) begin
					state<=2;
					out<=193;
				end
				if(in == 924) begin
					state<=2;
					out<=194;
				end
				if(in == 925) begin
					state<=2;
					out<=195;
				end
				if(in == 926) begin
					state<=2;
					out<=196;
				end
				if(in == 927) begin
					state<=2;
					out<=197;
				end
				if(in == 928) begin
					state<=2;
					out<=198;
				end
			end
			7: begin
				if(in == 0) begin
					state<=3;
					out<=199;
				end
				if(in == 1) begin
					state<=1;
					out<=200;
				end
				if(in == 2) begin
					state<=7;
					out<=201;
				end
				if(in == 3) begin
					state<=3;
					out<=202;
				end
				if(in == 4) begin
					state<=12;
					out<=203;
				end
				if(in == 5) begin
					state<=3;
					out<=204;
				end
				if(in == 6) begin
					state<=12;
					out<=205;
				end
				if(in == 7) begin
					state<=12;
					out<=206;
				end
				if(in == 8) begin
					state<=12;
					out<=207;
				end
				if(in == 9) begin
					state<=18;
					out<=208;
				end
				if(in == 10) begin
					state<=18;
					out<=209;
				end
				if(in == 11) begin
					state<=18;
					out<=210;
				end
				if(in == 12) begin
					state<=18;
					out<=211;
				end
				if(in == 13) begin
					state<=24;
					out<=212;
				end
				if(in == 14) begin
					state<=24;
					out<=213;
				end
				if(in == 15) begin
					state<=24;
					out<=214;
				end
				if(in == 16) begin
					state<=24;
					out<=215;
				end
				if(in == 17) begin
					state<=8;
					out<=216;
				end
				if(in == 18) begin
					state<=8;
					out<=217;
				end
				if(in == 19) begin
					state<=8;
					out<=218;
				end
				if(in == 20) begin
					state<=8;
					out<=219;
				end
				if(in == 21) begin
					state<=12;
					out<=220;
				end
				if(in == 22) begin
					state<=12;
					out<=221;
				end
				if(in == 23) begin
					state<=12;
					out<=222;
				end
				if(in == 24) begin
					state<=12;
					out<=223;
				end
				if(in == 25) begin
					state<=18;
					out<=224;
				end
				if(in == 26) begin
					state<=18;
					out<=225;
				end
				if(in == 27) begin
					state<=18;
					out<=226;
				end
				if(in == 28) begin
					state<=18;
					out<=227;
				end
				if(in == 29) begin
					state<=24;
					out<=228;
				end
				if(in == 30) begin
					state<=24;
					out<=229;
				end
				if(in == 31) begin
					state<=24;
					out<=230;
				end
				if(in == 32) begin
					state<=24;
					out<=231;
				end
				if(in == 33) begin
					state<=8;
					out<=232;
				end
				if(in == 34) begin
					state<=8;
					out<=233;
				end
				if(in == 35) begin
					state<=8;
					out<=234;
				end
				if(in == 36) begin
					state<=8;
					out<=235;
				end
				if(in == 37) begin
					state<=12;
					out<=236;
				end
				if(in == 38) begin
					state<=12;
					out<=237;
				end
				if(in == 39) begin
					state<=12;
					out<=238;
				end
				if(in == 40) begin
					state<=12;
					out<=239;
				end
				if(in == 41) begin
					state<=18;
					out<=240;
				end
				if(in == 42) begin
					state<=18;
					out<=241;
				end
				if(in == 43) begin
					state<=18;
					out<=242;
				end
				if(in == 44) begin
					state<=18;
					out<=243;
				end
				if(in == 45) begin
					state<=24;
					out<=244;
				end
				if(in == 46) begin
					state<=24;
					out<=245;
				end
				if(in == 47) begin
					state<=24;
					out<=246;
				end
				if(in == 48) begin
					state<=24;
					out<=247;
				end
				if(in == 49) begin
					state<=8;
					out<=248;
				end
				if(in == 50) begin
					state<=8;
					out<=249;
				end
				if(in == 51) begin
					state<=8;
					out<=250;
				end
				if(in == 52) begin
					state<=8;
					out<=251;
				end
				if(in == 53) begin
					state<=3;
					out<=252;
				end
				if(in == 54) begin
					state<=7;
					out<=253;
				end
				if(in == 55) begin
					state<=3;
					out<=254;
				end
				if(in == 56) begin
					state<=12;
					out<=255;
				end
				if(in == 57) begin
					state<=3;
					out<=0;
				end
				if(in == 58) begin
					state<=12;
					out<=1;
				end
				if(in == 59) begin
					state<=12;
					out<=2;
				end
				if(in == 60) begin
					state<=12;
					out<=3;
				end
				if(in == 61) begin
					state<=18;
					out<=4;
				end
				if(in == 62) begin
					state<=18;
					out<=5;
				end
				if(in == 63) begin
					state<=18;
					out<=6;
				end
				if(in == 64) begin
					state<=18;
					out<=7;
				end
				if(in == 65) begin
					state<=24;
					out<=8;
				end
				if(in == 66) begin
					state<=24;
					out<=9;
				end
				if(in == 67) begin
					state<=24;
					out<=10;
				end
				if(in == 68) begin
					state<=24;
					out<=11;
				end
				if(in == 69) begin
					state<=8;
					out<=12;
				end
				if(in == 70) begin
					state<=8;
					out<=13;
				end
				if(in == 71) begin
					state<=8;
					out<=14;
				end
				if(in == 72) begin
					state<=8;
					out<=15;
				end
				if(in == 73) begin
					state<=12;
					out<=16;
				end
				if(in == 74) begin
					state<=12;
					out<=17;
				end
				if(in == 75) begin
					state<=12;
					out<=18;
				end
				if(in == 76) begin
					state<=12;
					out<=19;
				end
				if(in == 77) begin
					state<=18;
					out<=20;
				end
				if(in == 78) begin
					state<=18;
					out<=21;
				end
				if(in == 79) begin
					state<=18;
					out<=22;
				end
				if(in == 80) begin
					state<=18;
					out<=23;
				end
				if(in == 81) begin
					state<=24;
					out<=24;
				end
				if(in == 82) begin
					state<=24;
					out<=25;
				end
				if(in == 83) begin
					state<=24;
					out<=26;
				end
				if(in == 84) begin
					state<=24;
					out<=27;
				end
				if(in == 85) begin
					state<=8;
					out<=28;
				end
				if(in == 86) begin
					state<=8;
					out<=29;
				end
				if(in == 87) begin
					state<=8;
					out<=30;
				end
				if(in == 88) begin
					state<=8;
					out<=31;
				end
				if(in == 89) begin
					state<=12;
					out<=32;
				end
				if(in == 90) begin
					state<=12;
					out<=33;
				end
				if(in == 91) begin
					state<=12;
					out<=34;
				end
				if(in == 92) begin
					state<=12;
					out<=35;
				end
				if(in == 93) begin
					state<=18;
					out<=36;
				end
				if(in == 94) begin
					state<=18;
					out<=37;
				end
				if(in == 95) begin
					state<=18;
					out<=38;
				end
				if(in == 96) begin
					state<=18;
					out<=39;
				end
				if(in == 97) begin
					state<=24;
					out<=40;
				end
				if(in == 98) begin
					state<=24;
					out<=41;
				end
				if(in == 99) begin
					state<=24;
					out<=42;
				end
				if(in == 100) begin
					state<=24;
					out<=43;
				end
				if(in == 101) begin
					state<=8;
					out<=44;
				end
				if(in == 102) begin
					state<=8;
					out<=45;
				end
				if(in == 103) begin
					state<=8;
					out<=46;
				end
				if(in == 104) begin
					state<=8;
					out<=47;
				end
				if(in == 105) begin
					state<=2;
					out<=48;
				end
				if(in == 106) begin
					state<=2;
					out<=49;
				end
				if(in == 107) begin
					state<=2;
					out<=50;
				end
				if(in == 108) begin
					state<=2;
					out<=51;
				end
				if(in == 109) begin
					state<=2;
					out<=52;
				end
				if(in == 110) begin
					state<=2;
					out<=53;
				end
				if(in == 111) begin
					state<=2;
					out<=54;
				end
				if(in == 112) begin
					state<=2;
					out<=55;
				end
				if(in == 113) begin
					state<=2;
					out<=56;
				end
				if(in == 114) begin
					state<=2;
					out<=57;
				end
				if(in == 115) begin
					state<=2;
					out<=58;
				end
				if(in == 116) begin
					state<=2;
					out<=59;
				end
				if(in == 117) begin
					state<=3;
					out<=60;
				end
				if(in == 118) begin
					state<=7;
					out<=61;
				end
				if(in == 119) begin
					state<=3;
					out<=62;
				end
				if(in == 120) begin
					state<=12;
					out<=63;
				end
				if(in == 121) begin
					state<=3;
					out<=64;
				end
				if(in == 122) begin
					state<=12;
					out<=65;
				end
				if(in == 123) begin
					state<=12;
					out<=66;
				end
				if(in == 124) begin
					state<=12;
					out<=67;
				end
				if(in == 125) begin
					state<=18;
					out<=68;
				end
				if(in == 126) begin
					state<=18;
					out<=69;
				end
				if(in == 127) begin
					state<=18;
					out<=70;
				end
				if(in == 128) begin
					state<=18;
					out<=71;
				end
				if(in == 129) begin
					state<=24;
					out<=72;
				end
				if(in == 130) begin
					state<=24;
					out<=73;
				end
				if(in == 131) begin
					state<=24;
					out<=74;
				end
				if(in == 132) begin
					state<=24;
					out<=75;
				end
				if(in == 133) begin
					state<=8;
					out<=76;
				end
				if(in == 134) begin
					state<=8;
					out<=77;
				end
				if(in == 135) begin
					state<=8;
					out<=78;
				end
				if(in == 136) begin
					state<=8;
					out<=79;
				end
				if(in == 137) begin
					state<=12;
					out<=80;
				end
				if(in == 138) begin
					state<=12;
					out<=81;
				end
				if(in == 139) begin
					state<=12;
					out<=82;
				end
				if(in == 140) begin
					state<=12;
					out<=83;
				end
				if(in == 141) begin
					state<=18;
					out<=84;
				end
				if(in == 142) begin
					state<=18;
					out<=85;
				end
				if(in == 143) begin
					state<=18;
					out<=86;
				end
				if(in == 144) begin
					state<=18;
					out<=87;
				end
				if(in == 145) begin
					state<=24;
					out<=88;
				end
				if(in == 146) begin
					state<=24;
					out<=89;
				end
				if(in == 147) begin
					state<=24;
					out<=90;
				end
				if(in == 148) begin
					state<=24;
					out<=91;
				end
				if(in == 149) begin
					state<=8;
					out<=92;
				end
				if(in == 150) begin
					state<=8;
					out<=93;
				end
				if(in == 151) begin
					state<=8;
					out<=94;
				end
				if(in == 152) begin
					state<=8;
					out<=95;
				end
				if(in == 153) begin
					state<=12;
					out<=96;
				end
				if(in == 154) begin
					state<=12;
					out<=97;
				end
				if(in == 155) begin
					state<=12;
					out<=98;
				end
				if(in == 156) begin
					state<=12;
					out<=99;
				end
				if(in == 157) begin
					state<=18;
					out<=100;
				end
				if(in == 158) begin
					state<=18;
					out<=101;
				end
				if(in == 159) begin
					state<=18;
					out<=102;
				end
				if(in == 160) begin
					state<=18;
					out<=103;
				end
				if(in == 161) begin
					state<=24;
					out<=104;
				end
				if(in == 162) begin
					state<=24;
					out<=105;
				end
				if(in == 163) begin
					state<=24;
					out<=106;
				end
				if(in == 164) begin
					state<=24;
					out<=107;
				end
				if(in == 165) begin
					state<=8;
					out<=108;
				end
				if(in == 166) begin
					state<=8;
					out<=109;
				end
				if(in == 167) begin
					state<=8;
					out<=110;
				end
				if(in == 168) begin
					state<=8;
					out<=111;
				end
				if(in == 169) begin
					state<=3;
					out<=112;
				end
				if(in == 170) begin
					state<=7;
					out<=113;
				end
				if(in == 171) begin
					state<=3;
					out<=114;
				end
				if(in == 172) begin
					state<=12;
					out<=115;
				end
				if(in == 173) begin
					state<=3;
					out<=116;
				end
				if(in == 174) begin
					state<=12;
					out<=117;
				end
				if(in == 175) begin
					state<=12;
					out<=118;
				end
				if(in == 176) begin
					state<=12;
					out<=119;
				end
				if(in == 177) begin
					state<=18;
					out<=120;
				end
				if(in == 178) begin
					state<=18;
					out<=121;
				end
				if(in == 179) begin
					state<=18;
					out<=122;
				end
				if(in == 180) begin
					state<=18;
					out<=123;
				end
				if(in == 181) begin
					state<=24;
					out<=124;
				end
				if(in == 182) begin
					state<=24;
					out<=125;
				end
				if(in == 183) begin
					state<=24;
					out<=126;
				end
				if(in == 184) begin
					state<=24;
					out<=127;
				end
				if(in == 185) begin
					state<=8;
					out<=128;
				end
				if(in == 186) begin
					state<=8;
					out<=129;
				end
				if(in == 187) begin
					state<=8;
					out<=130;
				end
				if(in == 188) begin
					state<=8;
					out<=131;
				end
				if(in == 189) begin
					state<=12;
					out<=132;
				end
				if(in == 190) begin
					state<=12;
					out<=133;
				end
				if(in == 191) begin
					state<=12;
					out<=134;
				end
				if(in == 192) begin
					state<=12;
					out<=135;
				end
				if(in == 193) begin
					state<=18;
					out<=136;
				end
				if(in == 194) begin
					state<=18;
					out<=137;
				end
				if(in == 195) begin
					state<=18;
					out<=138;
				end
				if(in == 196) begin
					state<=18;
					out<=139;
				end
				if(in == 197) begin
					state<=24;
					out<=140;
				end
				if(in == 198) begin
					state<=24;
					out<=141;
				end
				if(in == 199) begin
					state<=24;
					out<=142;
				end
				if(in == 200) begin
					state<=24;
					out<=143;
				end
				if(in == 201) begin
					state<=8;
					out<=144;
				end
				if(in == 202) begin
					state<=8;
					out<=145;
				end
				if(in == 203) begin
					state<=8;
					out<=146;
				end
				if(in == 204) begin
					state<=8;
					out<=147;
				end
				if(in == 205) begin
					state<=12;
					out<=148;
				end
				if(in == 206) begin
					state<=12;
					out<=149;
				end
				if(in == 207) begin
					state<=12;
					out<=150;
				end
				if(in == 208) begin
					state<=12;
					out<=151;
				end
				if(in == 209) begin
					state<=18;
					out<=152;
				end
				if(in == 210) begin
					state<=18;
					out<=153;
				end
				if(in == 211) begin
					state<=18;
					out<=154;
				end
				if(in == 212) begin
					state<=18;
					out<=155;
				end
				if(in == 213) begin
					state<=24;
					out<=156;
				end
				if(in == 214) begin
					state<=24;
					out<=157;
				end
				if(in == 215) begin
					state<=24;
					out<=158;
				end
				if(in == 216) begin
					state<=24;
					out<=159;
				end
				if(in == 217) begin
					state<=8;
					out<=160;
				end
				if(in == 218) begin
					state<=8;
					out<=161;
				end
				if(in == 219) begin
					state<=8;
					out<=162;
				end
				if(in == 220) begin
					state<=8;
					out<=163;
				end
				if(in == 221) begin
					state<=2;
					out<=164;
				end
				if(in == 222) begin
					state<=2;
					out<=165;
				end
				if(in == 223) begin
					state<=2;
					out<=166;
				end
				if(in == 224) begin
					state<=2;
					out<=167;
				end
				if(in == 225) begin
					state<=2;
					out<=168;
				end
				if(in == 226) begin
					state<=2;
					out<=169;
				end
				if(in == 227) begin
					state<=2;
					out<=170;
				end
				if(in == 228) begin
					state<=2;
					out<=171;
				end
				if(in == 229) begin
					state<=2;
					out<=172;
				end
				if(in == 230) begin
					state<=2;
					out<=173;
				end
				if(in == 231) begin
					state<=2;
					out<=174;
				end
				if(in == 232) begin
					state<=2;
					out<=175;
				end
				if(in == 233) begin
					state<=3;
					out<=176;
				end
				if(in == 234) begin
					state<=7;
					out<=177;
				end
				if(in == 235) begin
					state<=3;
					out<=178;
				end
				if(in == 236) begin
					state<=12;
					out<=179;
				end
				if(in == 237) begin
					state<=3;
					out<=180;
				end
				if(in == 238) begin
					state<=12;
					out<=181;
				end
				if(in == 239) begin
					state<=12;
					out<=182;
				end
				if(in == 240) begin
					state<=12;
					out<=183;
				end
				if(in == 241) begin
					state<=18;
					out<=184;
				end
				if(in == 242) begin
					state<=18;
					out<=185;
				end
				if(in == 243) begin
					state<=18;
					out<=186;
				end
				if(in == 244) begin
					state<=18;
					out<=187;
				end
				if(in == 245) begin
					state<=24;
					out<=188;
				end
				if(in == 246) begin
					state<=24;
					out<=189;
				end
				if(in == 247) begin
					state<=24;
					out<=190;
				end
				if(in == 248) begin
					state<=24;
					out<=191;
				end
				if(in == 249) begin
					state<=8;
					out<=192;
				end
				if(in == 250) begin
					state<=8;
					out<=193;
				end
				if(in == 251) begin
					state<=8;
					out<=194;
				end
				if(in == 252) begin
					state<=8;
					out<=195;
				end
				if(in == 253) begin
					state<=12;
					out<=196;
				end
				if(in == 254) begin
					state<=12;
					out<=197;
				end
				if(in == 255) begin
					state<=12;
					out<=198;
				end
				if(in == 256) begin
					state<=12;
					out<=199;
				end
				if(in == 257) begin
					state<=18;
					out<=200;
				end
				if(in == 258) begin
					state<=18;
					out<=201;
				end
				if(in == 259) begin
					state<=18;
					out<=202;
				end
				if(in == 260) begin
					state<=18;
					out<=203;
				end
				if(in == 261) begin
					state<=24;
					out<=204;
				end
				if(in == 262) begin
					state<=24;
					out<=205;
				end
				if(in == 263) begin
					state<=24;
					out<=206;
				end
				if(in == 264) begin
					state<=24;
					out<=207;
				end
				if(in == 265) begin
					state<=8;
					out<=208;
				end
				if(in == 266) begin
					state<=8;
					out<=209;
				end
				if(in == 267) begin
					state<=8;
					out<=210;
				end
				if(in == 268) begin
					state<=8;
					out<=211;
				end
				if(in == 269) begin
					state<=12;
					out<=212;
				end
				if(in == 270) begin
					state<=12;
					out<=213;
				end
				if(in == 271) begin
					state<=12;
					out<=214;
				end
				if(in == 272) begin
					state<=12;
					out<=215;
				end
				if(in == 273) begin
					state<=18;
					out<=216;
				end
				if(in == 274) begin
					state<=18;
					out<=217;
				end
				if(in == 275) begin
					state<=18;
					out<=218;
				end
				if(in == 276) begin
					state<=18;
					out<=219;
				end
				if(in == 277) begin
					state<=24;
					out<=220;
				end
				if(in == 278) begin
					state<=24;
					out<=221;
				end
				if(in == 279) begin
					state<=24;
					out<=222;
				end
				if(in == 280) begin
					state<=24;
					out<=223;
				end
				if(in == 281) begin
					state<=8;
					out<=224;
				end
				if(in == 282) begin
					state<=8;
					out<=225;
				end
				if(in == 283) begin
					state<=8;
					out<=226;
				end
				if(in == 284) begin
					state<=8;
					out<=227;
				end
				if(in == 285) begin
					state<=3;
					out<=228;
				end
				if(in == 286) begin
					state<=7;
					out<=229;
				end
				if(in == 287) begin
					state<=3;
					out<=230;
				end
				if(in == 288) begin
					state<=12;
					out<=231;
				end
				if(in == 289) begin
					state<=3;
					out<=232;
				end
				if(in == 290) begin
					state<=12;
					out<=233;
				end
				if(in == 291) begin
					state<=12;
					out<=234;
				end
				if(in == 292) begin
					state<=12;
					out<=235;
				end
				if(in == 293) begin
					state<=18;
					out<=236;
				end
				if(in == 294) begin
					state<=18;
					out<=237;
				end
				if(in == 295) begin
					state<=18;
					out<=238;
				end
				if(in == 296) begin
					state<=18;
					out<=239;
				end
				if(in == 297) begin
					state<=24;
					out<=240;
				end
				if(in == 298) begin
					state<=24;
					out<=241;
				end
				if(in == 299) begin
					state<=24;
					out<=242;
				end
				if(in == 300) begin
					state<=24;
					out<=243;
				end
				if(in == 301) begin
					state<=8;
					out<=244;
				end
				if(in == 302) begin
					state<=8;
					out<=245;
				end
				if(in == 303) begin
					state<=8;
					out<=246;
				end
				if(in == 304) begin
					state<=8;
					out<=247;
				end
				if(in == 305) begin
					state<=12;
					out<=248;
				end
				if(in == 306) begin
					state<=12;
					out<=249;
				end
				if(in == 307) begin
					state<=12;
					out<=250;
				end
				if(in == 308) begin
					state<=12;
					out<=251;
				end
				if(in == 309) begin
					state<=18;
					out<=252;
				end
				if(in == 310) begin
					state<=18;
					out<=253;
				end
				if(in == 311) begin
					state<=18;
					out<=254;
				end
				if(in == 312) begin
					state<=18;
					out<=255;
				end
				if(in == 313) begin
					state<=24;
					out<=0;
				end
				if(in == 314) begin
					state<=24;
					out<=1;
				end
				if(in == 315) begin
					state<=24;
					out<=2;
				end
				if(in == 316) begin
					state<=24;
					out<=3;
				end
				if(in == 317) begin
					state<=8;
					out<=4;
				end
				if(in == 318) begin
					state<=8;
					out<=5;
				end
				if(in == 319) begin
					state<=8;
					out<=6;
				end
				if(in == 320) begin
					state<=8;
					out<=7;
				end
				if(in == 321) begin
					state<=12;
					out<=8;
				end
				if(in == 322) begin
					state<=12;
					out<=9;
				end
				if(in == 323) begin
					state<=12;
					out<=10;
				end
				if(in == 324) begin
					state<=12;
					out<=11;
				end
				if(in == 325) begin
					state<=18;
					out<=12;
				end
				if(in == 326) begin
					state<=18;
					out<=13;
				end
				if(in == 327) begin
					state<=18;
					out<=14;
				end
				if(in == 328) begin
					state<=18;
					out<=15;
				end
				if(in == 329) begin
					state<=24;
					out<=16;
				end
				if(in == 330) begin
					state<=24;
					out<=17;
				end
				if(in == 331) begin
					state<=24;
					out<=18;
				end
				if(in == 332) begin
					state<=24;
					out<=19;
				end
				if(in == 333) begin
					state<=8;
					out<=20;
				end
				if(in == 334) begin
					state<=8;
					out<=21;
				end
				if(in == 335) begin
					state<=8;
					out<=22;
				end
				if(in == 336) begin
					state<=8;
					out<=23;
				end
				if(in == 337) begin
					state<=2;
					out<=24;
				end
				if(in == 338) begin
					state<=2;
					out<=25;
				end
				if(in == 339) begin
					state<=2;
					out<=26;
				end
				if(in == 340) begin
					state<=2;
					out<=27;
				end
				if(in == 341) begin
					state<=2;
					out<=28;
				end
				if(in == 342) begin
					state<=2;
					out<=29;
				end
				if(in == 343) begin
					state<=2;
					out<=30;
				end
				if(in == 344) begin
					state<=2;
					out<=31;
				end
				if(in == 345) begin
					state<=2;
					out<=32;
				end
				if(in == 346) begin
					state<=2;
					out<=33;
				end
				if(in == 347) begin
					state<=2;
					out<=34;
				end
				if(in == 348) begin
					state<=2;
					out<=35;
				end
				if(in == 349) begin
					state<=3;
					out<=36;
				end
				if(in == 350) begin
					state<=7;
					out<=37;
				end
				if(in == 351) begin
					state<=3;
					out<=38;
				end
				if(in == 352) begin
					state<=12;
					out<=39;
				end
				if(in == 353) begin
					state<=3;
					out<=40;
				end
				if(in == 354) begin
					state<=12;
					out<=41;
				end
				if(in == 355) begin
					state<=12;
					out<=42;
				end
				if(in == 356) begin
					state<=12;
					out<=43;
				end
				if(in == 357) begin
					state<=18;
					out<=44;
				end
				if(in == 358) begin
					state<=18;
					out<=45;
				end
				if(in == 359) begin
					state<=18;
					out<=46;
				end
				if(in == 360) begin
					state<=18;
					out<=47;
				end
				if(in == 361) begin
					state<=24;
					out<=48;
				end
				if(in == 362) begin
					state<=24;
					out<=49;
				end
				if(in == 363) begin
					state<=24;
					out<=50;
				end
				if(in == 364) begin
					state<=24;
					out<=51;
				end
				if(in == 365) begin
					state<=8;
					out<=52;
				end
				if(in == 366) begin
					state<=8;
					out<=53;
				end
				if(in == 367) begin
					state<=8;
					out<=54;
				end
				if(in == 368) begin
					state<=8;
					out<=55;
				end
				if(in == 369) begin
					state<=12;
					out<=56;
				end
				if(in == 370) begin
					state<=12;
					out<=57;
				end
				if(in == 371) begin
					state<=12;
					out<=58;
				end
				if(in == 372) begin
					state<=12;
					out<=59;
				end
				if(in == 373) begin
					state<=18;
					out<=60;
				end
				if(in == 374) begin
					state<=18;
					out<=61;
				end
				if(in == 375) begin
					state<=18;
					out<=62;
				end
				if(in == 376) begin
					state<=18;
					out<=63;
				end
				if(in == 377) begin
					state<=24;
					out<=64;
				end
				if(in == 378) begin
					state<=24;
					out<=65;
				end
				if(in == 379) begin
					state<=24;
					out<=66;
				end
				if(in == 380) begin
					state<=24;
					out<=67;
				end
				if(in == 381) begin
					state<=8;
					out<=68;
				end
				if(in == 382) begin
					state<=8;
					out<=69;
				end
				if(in == 383) begin
					state<=8;
					out<=70;
				end
				if(in == 384) begin
					state<=8;
					out<=71;
				end
				if(in == 385) begin
					state<=12;
					out<=72;
				end
				if(in == 386) begin
					state<=12;
					out<=73;
				end
				if(in == 387) begin
					state<=12;
					out<=74;
				end
				if(in == 388) begin
					state<=12;
					out<=75;
				end
				if(in == 389) begin
					state<=18;
					out<=76;
				end
				if(in == 390) begin
					state<=18;
					out<=77;
				end
				if(in == 391) begin
					state<=18;
					out<=78;
				end
				if(in == 392) begin
					state<=18;
					out<=79;
				end
				if(in == 393) begin
					state<=24;
					out<=80;
				end
				if(in == 394) begin
					state<=24;
					out<=81;
				end
				if(in == 395) begin
					state<=24;
					out<=82;
				end
				if(in == 396) begin
					state<=24;
					out<=83;
				end
				if(in == 397) begin
					state<=8;
					out<=84;
				end
				if(in == 398) begin
					state<=8;
					out<=85;
				end
				if(in == 399) begin
					state<=8;
					out<=86;
				end
				if(in == 400) begin
					state<=8;
					out<=87;
				end
				if(in == 401) begin
					state<=3;
					out<=88;
				end
				if(in == 402) begin
					state<=7;
					out<=89;
				end
				if(in == 403) begin
					state<=3;
					out<=90;
				end
				if(in == 404) begin
					state<=12;
					out<=91;
				end
				if(in == 405) begin
					state<=3;
					out<=92;
				end
				if(in == 406) begin
					state<=12;
					out<=93;
				end
				if(in == 407) begin
					state<=12;
					out<=94;
				end
				if(in == 408) begin
					state<=12;
					out<=95;
				end
				if(in == 409) begin
					state<=18;
					out<=96;
				end
				if(in == 410) begin
					state<=18;
					out<=97;
				end
				if(in == 411) begin
					state<=18;
					out<=98;
				end
				if(in == 412) begin
					state<=18;
					out<=99;
				end
				if(in == 413) begin
					state<=24;
					out<=100;
				end
				if(in == 414) begin
					state<=24;
					out<=101;
				end
				if(in == 415) begin
					state<=24;
					out<=102;
				end
				if(in == 416) begin
					state<=24;
					out<=103;
				end
				if(in == 417) begin
					state<=8;
					out<=104;
				end
				if(in == 418) begin
					state<=8;
					out<=105;
				end
				if(in == 419) begin
					state<=8;
					out<=106;
				end
				if(in == 420) begin
					state<=8;
					out<=107;
				end
				if(in == 421) begin
					state<=12;
					out<=108;
				end
				if(in == 422) begin
					state<=12;
					out<=109;
				end
				if(in == 423) begin
					state<=12;
					out<=110;
				end
				if(in == 424) begin
					state<=12;
					out<=111;
				end
				if(in == 425) begin
					state<=18;
					out<=112;
				end
				if(in == 426) begin
					state<=18;
					out<=113;
				end
				if(in == 427) begin
					state<=18;
					out<=114;
				end
				if(in == 428) begin
					state<=18;
					out<=115;
				end
				if(in == 429) begin
					state<=24;
					out<=116;
				end
				if(in == 430) begin
					state<=24;
					out<=117;
				end
				if(in == 431) begin
					state<=24;
					out<=118;
				end
				if(in == 432) begin
					state<=24;
					out<=119;
				end
				if(in == 433) begin
					state<=8;
					out<=120;
				end
				if(in == 434) begin
					state<=8;
					out<=121;
				end
				if(in == 435) begin
					state<=8;
					out<=122;
				end
				if(in == 436) begin
					state<=8;
					out<=123;
				end
				if(in == 437) begin
					state<=12;
					out<=124;
				end
				if(in == 438) begin
					state<=12;
					out<=125;
				end
				if(in == 439) begin
					state<=12;
					out<=126;
				end
				if(in == 440) begin
					state<=12;
					out<=127;
				end
				if(in == 441) begin
					state<=18;
					out<=128;
				end
				if(in == 442) begin
					state<=18;
					out<=129;
				end
				if(in == 443) begin
					state<=18;
					out<=130;
				end
				if(in == 444) begin
					state<=18;
					out<=131;
				end
				if(in == 445) begin
					state<=24;
					out<=132;
				end
				if(in == 446) begin
					state<=24;
					out<=133;
				end
				if(in == 447) begin
					state<=24;
					out<=134;
				end
				if(in == 448) begin
					state<=24;
					out<=135;
				end
				if(in == 449) begin
					state<=8;
					out<=136;
				end
				if(in == 450) begin
					state<=8;
					out<=137;
				end
				if(in == 451) begin
					state<=8;
					out<=138;
				end
				if(in == 452) begin
					state<=8;
					out<=139;
				end
				if(in == 453) begin
					state<=2;
					out<=140;
				end
				if(in == 454) begin
					state<=2;
					out<=141;
				end
				if(in == 455) begin
					state<=2;
					out<=142;
				end
				if(in == 456) begin
					state<=2;
					out<=143;
				end
				if(in == 457) begin
					state<=2;
					out<=144;
				end
				if(in == 458) begin
					state<=2;
					out<=145;
				end
				if(in == 459) begin
					state<=2;
					out<=146;
				end
				if(in == 460) begin
					state<=2;
					out<=147;
				end
				if(in == 461) begin
					state<=2;
					out<=148;
				end
				if(in == 462) begin
					state<=2;
					out<=149;
				end
				if(in == 463) begin
					state<=2;
					out<=150;
				end
				if(in == 464) begin
					state<=2;
					out<=151;
				end
				if(in == 465) begin
					state<=3;
					out<=152;
				end
				if(in == 466) begin
					state<=7;
					out<=153;
				end
				if(in == 467) begin
					state<=3;
					out<=154;
				end
				if(in == 468) begin
					state<=12;
					out<=155;
				end
				if(in == 469) begin
					state<=3;
					out<=156;
				end
				if(in == 470) begin
					state<=12;
					out<=157;
				end
				if(in == 471) begin
					state<=12;
					out<=158;
				end
				if(in == 472) begin
					state<=12;
					out<=159;
				end
				if(in == 473) begin
					state<=18;
					out<=160;
				end
				if(in == 474) begin
					state<=18;
					out<=161;
				end
				if(in == 475) begin
					state<=18;
					out<=162;
				end
				if(in == 476) begin
					state<=18;
					out<=163;
				end
				if(in == 477) begin
					state<=24;
					out<=164;
				end
				if(in == 478) begin
					state<=24;
					out<=165;
				end
				if(in == 479) begin
					state<=24;
					out<=166;
				end
				if(in == 480) begin
					state<=24;
					out<=167;
				end
				if(in == 481) begin
					state<=8;
					out<=168;
				end
				if(in == 482) begin
					state<=8;
					out<=169;
				end
				if(in == 483) begin
					state<=8;
					out<=170;
				end
				if(in == 484) begin
					state<=8;
					out<=171;
				end
				if(in == 485) begin
					state<=12;
					out<=172;
				end
				if(in == 486) begin
					state<=12;
					out<=173;
				end
				if(in == 487) begin
					state<=12;
					out<=174;
				end
				if(in == 488) begin
					state<=12;
					out<=175;
				end
				if(in == 489) begin
					state<=18;
					out<=176;
				end
				if(in == 490) begin
					state<=18;
					out<=177;
				end
				if(in == 491) begin
					state<=18;
					out<=178;
				end
				if(in == 492) begin
					state<=18;
					out<=179;
				end
				if(in == 493) begin
					state<=24;
					out<=180;
				end
				if(in == 494) begin
					state<=24;
					out<=181;
				end
				if(in == 495) begin
					state<=24;
					out<=182;
				end
				if(in == 496) begin
					state<=24;
					out<=183;
				end
				if(in == 497) begin
					state<=8;
					out<=184;
				end
				if(in == 498) begin
					state<=8;
					out<=185;
				end
				if(in == 499) begin
					state<=8;
					out<=186;
				end
				if(in == 500) begin
					state<=8;
					out<=187;
				end
				if(in == 501) begin
					state<=12;
					out<=188;
				end
				if(in == 502) begin
					state<=12;
					out<=189;
				end
				if(in == 503) begin
					state<=12;
					out<=190;
				end
				if(in == 504) begin
					state<=12;
					out<=191;
				end
				if(in == 505) begin
					state<=18;
					out<=192;
				end
				if(in == 506) begin
					state<=18;
					out<=193;
				end
				if(in == 507) begin
					state<=18;
					out<=194;
				end
				if(in == 508) begin
					state<=18;
					out<=195;
				end
				if(in == 509) begin
					state<=24;
					out<=196;
				end
				if(in == 510) begin
					state<=24;
					out<=197;
				end
				if(in == 511) begin
					state<=24;
					out<=198;
				end
				if(in == 512) begin
					state<=24;
					out<=199;
				end
				if(in == 513) begin
					state<=8;
					out<=200;
				end
				if(in == 514) begin
					state<=8;
					out<=201;
				end
				if(in == 515) begin
					state<=8;
					out<=202;
				end
				if(in == 516) begin
					state<=8;
					out<=203;
				end
				if(in == 517) begin
					state<=3;
					out<=204;
				end
				if(in == 518) begin
					state<=7;
					out<=205;
				end
				if(in == 519) begin
					state<=3;
					out<=206;
				end
				if(in == 520) begin
					state<=12;
					out<=207;
				end
				if(in == 521) begin
					state<=3;
					out<=208;
				end
				if(in == 522) begin
					state<=12;
					out<=209;
				end
				if(in == 523) begin
					state<=12;
					out<=210;
				end
				if(in == 524) begin
					state<=12;
					out<=211;
				end
				if(in == 525) begin
					state<=18;
					out<=212;
				end
				if(in == 526) begin
					state<=18;
					out<=213;
				end
				if(in == 527) begin
					state<=18;
					out<=214;
				end
				if(in == 528) begin
					state<=18;
					out<=215;
				end
				if(in == 529) begin
					state<=24;
					out<=216;
				end
				if(in == 530) begin
					state<=24;
					out<=217;
				end
				if(in == 531) begin
					state<=24;
					out<=218;
				end
				if(in == 532) begin
					state<=24;
					out<=219;
				end
				if(in == 533) begin
					state<=8;
					out<=220;
				end
				if(in == 534) begin
					state<=8;
					out<=221;
				end
				if(in == 535) begin
					state<=8;
					out<=222;
				end
				if(in == 536) begin
					state<=8;
					out<=223;
				end
				if(in == 537) begin
					state<=12;
					out<=224;
				end
				if(in == 538) begin
					state<=12;
					out<=225;
				end
				if(in == 539) begin
					state<=12;
					out<=226;
				end
				if(in == 540) begin
					state<=12;
					out<=227;
				end
				if(in == 541) begin
					state<=18;
					out<=228;
				end
				if(in == 542) begin
					state<=18;
					out<=229;
				end
				if(in == 543) begin
					state<=18;
					out<=230;
				end
				if(in == 544) begin
					state<=18;
					out<=231;
				end
				if(in == 545) begin
					state<=24;
					out<=232;
				end
				if(in == 546) begin
					state<=24;
					out<=233;
				end
				if(in == 547) begin
					state<=24;
					out<=234;
				end
				if(in == 548) begin
					state<=24;
					out<=235;
				end
				if(in == 549) begin
					state<=8;
					out<=236;
				end
				if(in == 550) begin
					state<=8;
					out<=237;
				end
				if(in == 551) begin
					state<=8;
					out<=238;
				end
				if(in == 552) begin
					state<=8;
					out<=239;
				end
				if(in == 553) begin
					state<=12;
					out<=240;
				end
				if(in == 554) begin
					state<=12;
					out<=241;
				end
				if(in == 555) begin
					state<=12;
					out<=242;
				end
				if(in == 556) begin
					state<=12;
					out<=243;
				end
				if(in == 557) begin
					state<=18;
					out<=244;
				end
				if(in == 558) begin
					state<=18;
					out<=245;
				end
				if(in == 559) begin
					state<=18;
					out<=246;
				end
				if(in == 560) begin
					state<=18;
					out<=247;
				end
				if(in == 561) begin
					state<=24;
					out<=248;
				end
				if(in == 562) begin
					state<=24;
					out<=249;
				end
				if(in == 563) begin
					state<=24;
					out<=250;
				end
				if(in == 564) begin
					state<=24;
					out<=251;
				end
				if(in == 565) begin
					state<=8;
					out<=252;
				end
				if(in == 566) begin
					state<=8;
					out<=253;
				end
				if(in == 567) begin
					state<=8;
					out<=254;
				end
				if(in == 568) begin
					state<=8;
					out<=255;
				end
				if(in == 569) begin
					state<=2;
					out<=0;
				end
				if(in == 570) begin
					state<=2;
					out<=1;
				end
				if(in == 571) begin
					state<=2;
					out<=2;
				end
				if(in == 572) begin
					state<=2;
					out<=3;
				end
				if(in == 573) begin
					state<=2;
					out<=4;
				end
				if(in == 574) begin
					state<=2;
					out<=5;
				end
				if(in == 575) begin
					state<=2;
					out<=6;
				end
				if(in == 576) begin
					state<=2;
					out<=7;
				end
				if(in == 577) begin
					state<=2;
					out<=8;
				end
				if(in == 578) begin
					state<=2;
					out<=9;
				end
				if(in == 579) begin
					state<=2;
					out<=10;
				end
				if(in == 580) begin
					state<=2;
					out<=11;
				end
				if(in == 581) begin
					state<=3;
					out<=12;
				end
				if(in == 582) begin
					state<=7;
					out<=13;
				end
				if(in == 583) begin
					state<=3;
					out<=14;
				end
				if(in == 584) begin
					state<=12;
					out<=15;
				end
				if(in == 585) begin
					state<=3;
					out<=16;
				end
				if(in == 586) begin
					state<=12;
					out<=17;
				end
				if(in == 587) begin
					state<=12;
					out<=18;
				end
				if(in == 588) begin
					state<=12;
					out<=19;
				end
				if(in == 589) begin
					state<=18;
					out<=20;
				end
				if(in == 590) begin
					state<=18;
					out<=21;
				end
				if(in == 591) begin
					state<=18;
					out<=22;
				end
				if(in == 592) begin
					state<=18;
					out<=23;
				end
				if(in == 593) begin
					state<=24;
					out<=24;
				end
				if(in == 594) begin
					state<=24;
					out<=25;
				end
				if(in == 595) begin
					state<=24;
					out<=26;
				end
				if(in == 596) begin
					state<=24;
					out<=27;
				end
				if(in == 597) begin
					state<=8;
					out<=28;
				end
				if(in == 598) begin
					state<=8;
					out<=29;
				end
				if(in == 599) begin
					state<=8;
					out<=30;
				end
				if(in == 600) begin
					state<=8;
					out<=31;
				end
				if(in == 601) begin
					state<=12;
					out<=32;
				end
				if(in == 602) begin
					state<=12;
					out<=33;
				end
				if(in == 603) begin
					state<=12;
					out<=34;
				end
				if(in == 604) begin
					state<=12;
					out<=35;
				end
				if(in == 605) begin
					state<=18;
					out<=36;
				end
				if(in == 606) begin
					state<=18;
					out<=37;
				end
				if(in == 607) begin
					state<=18;
					out<=38;
				end
				if(in == 608) begin
					state<=18;
					out<=39;
				end
				if(in == 609) begin
					state<=24;
					out<=40;
				end
				if(in == 610) begin
					state<=24;
					out<=41;
				end
				if(in == 611) begin
					state<=24;
					out<=42;
				end
				if(in == 612) begin
					state<=24;
					out<=43;
				end
				if(in == 613) begin
					state<=8;
					out<=44;
				end
				if(in == 614) begin
					state<=8;
					out<=45;
				end
				if(in == 615) begin
					state<=8;
					out<=46;
				end
				if(in == 616) begin
					state<=8;
					out<=47;
				end
				if(in == 617) begin
					state<=12;
					out<=48;
				end
				if(in == 618) begin
					state<=12;
					out<=49;
				end
				if(in == 619) begin
					state<=12;
					out<=50;
				end
				if(in == 620) begin
					state<=12;
					out<=51;
				end
				if(in == 621) begin
					state<=18;
					out<=52;
				end
				if(in == 622) begin
					state<=18;
					out<=53;
				end
				if(in == 623) begin
					state<=18;
					out<=54;
				end
				if(in == 624) begin
					state<=18;
					out<=55;
				end
				if(in == 625) begin
					state<=24;
					out<=56;
				end
				if(in == 626) begin
					state<=24;
					out<=57;
				end
				if(in == 627) begin
					state<=24;
					out<=58;
				end
				if(in == 628) begin
					state<=24;
					out<=59;
				end
				if(in == 629) begin
					state<=8;
					out<=60;
				end
				if(in == 630) begin
					state<=8;
					out<=61;
				end
				if(in == 631) begin
					state<=8;
					out<=62;
				end
				if(in == 632) begin
					state<=8;
					out<=63;
				end
				if(in == 633) begin
					state<=3;
					out<=64;
				end
				if(in == 634) begin
					state<=7;
					out<=65;
				end
				if(in == 635) begin
					state<=3;
					out<=66;
				end
				if(in == 636) begin
					state<=12;
					out<=67;
				end
				if(in == 637) begin
					state<=3;
					out<=68;
				end
				if(in == 638) begin
					state<=12;
					out<=69;
				end
				if(in == 639) begin
					state<=12;
					out<=70;
				end
				if(in == 640) begin
					state<=12;
					out<=71;
				end
				if(in == 641) begin
					state<=18;
					out<=72;
				end
				if(in == 642) begin
					state<=18;
					out<=73;
				end
				if(in == 643) begin
					state<=18;
					out<=74;
				end
				if(in == 644) begin
					state<=18;
					out<=75;
				end
				if(in == 645) begin
					state<=24;
					out<=76;
				end
				if(in == 646) begin
					state<=24;
					out<=77;
				end
				if(in == 647) begin
					state<=24;
					out<=78;
				end
				if(in == 648) begin
					state<=24;
					out<=79;
				end
				if(in == 649) begin
					state<=8;
					out<=80;
				end
				if(in == 650) begin
					state<=8;
					out<=81;
				end
				if(in == 651) begin
					state<=8;
					out<=82;
				end
				if(in == 652) begin
					state<=8;
					out<=83;
				end
				if(in == 653) begin
					state<=12;
					out<=84;
				end
				if(in == 654) begin
					state<=12;
					out<=85;
				end
				if(in == 655) begin
					state<=12;
					out<=86;
				end
				if(in == 656) begin
					state<=12;
					out<=87;
				end
				if(in == 657) begin
					state<=18;
					out<=88;
				end
				if(in == 658) begin
					state<=18;
					out<=89;
				end
				if(in == 659) begin
					state<=18;
					out<=90;
				end
				if(in == 660) begin
					state<=18;
					out<=91;
				end
				if(in == 661) begin
					state<=24;
					out<=92;
				end
				if(in == 662) begin
					state<=24;
					out<=93;
				end
				if(in == 663) begin
					state<=24;
					out<=94;
				end
				if(in == 664) begin
					state<=24;
					out<=95;
				end
				if(in == 665) begin
					state<=8;
					out<=96;
				end
				if(in == 666) begin
					state<=8;
					out<=97;
				end
				if(in == 667) begin
					state<=8;
					out<=98;
				end
				if(in == 668) begin
					state<=8;
					out<=99;
				end
				if(in == 669) begin
					state<=12;
					out<=100;
				end
				if(in == 670) begin
					state<=12;
					out<=101;
				end
				if(in == 671) begin
					state<=12;
					out<=102;
				end
				if(in == 672) begin
					state<=12;
					out<=103;
				end
				if(in == 673) begin
					state<=18;
					out<=104;
				end
				if(in == 674) begin
					state<=18;
					out<=105;
				end
				if(in == 675) begin
					state<=18;
					out<=106;
				end
				if(in == 676) begin
					state<=18;
					out<=107;
				end
				if(in == 677) begin
					state<=24;
					out<=108;
				end
				if(in == 678) begin
					state<=24;
					out<=109;
				end
				if(in == 679) begin
					state<=24;
					out<=110;
				end
				if(in == 680) begin
					state<=24;
					out<=111;
				end
				if(in == 681) begin
					state<=8;
					out<=112;
				end
				if(in == 682) begin
					state<=8;
					out<=113;
				end
				if(in == 683) begin
					state<=8;
					out<=114;
				end
				if(in == 684) begin
					state<=8;
					out<=115;
				end
				if(in == 685) begin
					state<=2;
					out<=116;
				end
				if(in == 686) begin
					state<=2;
					out<=117;
				end
				if(in == 687) begin
					state<=2;
					out<=118;
				end
				if(in == 688) begin
					state<=2;
					out<=119;
				end
				if(in == 689) begin
					state<=2;
					out<=120;
				end
				if(in == 690) begin
					state<=2;
					out<=121;
				end
				if(in == 691) begin
					state<=2;
					out<=122;
				end
				if(in == 692) begin
					state<=2;
					out<=123;
				end
				if(in == 693) begin
					state<=2;
					out<=124;
				end
				if(in == 694) begin
					state<=2;
					out<=125;
				end
				if(in == 695) begin
					state<=2;
					out<=126;
				end
				if(in == 696) begin
					state<=2;
					out<=127;
				end
				if(in == 697) begin
					state<=3;
					out<=128;
				end
				if(in == 698) begin
					state<=7;
					out<=129;
				end
				if(in == 699) begin
					state<=3;
					out<=130;
				end
				if(in == 700) begin
					state<=12;
					out<=131;
				end
				if(in == 701) begin
					state<=3;
					out<=132;
				end
				if(in == 702) begin
					state<=12;
					out<=133;
				end
				if(in == 703) begin
					state<=12;
					out<=134;
				end
				if(in == 704) begin
					state<=12;
					out<=135;
				end
				if(in == 705) begin
					state<=18;
					out<=136;
				end
				if(in == 706) begin
					state<=18;
					out<=137;
				end
				if(in == 707) begin
					state<=18;
					out<=138;
				end
				if(in == 708) begin
					state<=18;
					out<=139;
				end
				if(in == 709) begin
					state<=24;
					out<=140;
				end
				if(in == 710) begin
					state<=24;
					out<=141;
				end
				if(in == 711) begin
					state<=24;
					out<=142;
				end
				if(in == 712) begin
					state<=24;
					out<=143;
				end
				if(in == 713) begin
					state<=8;
					out<=144;
				end
				if(in == 714) begin
					state<=8;
					out<=145;
				end
				if(in == 715) begin
					state<=8;
					out<=146;
				end
				if(in == 716) begin
					state<=8;
					out<=147;
				end
				if(in == 717) begin
					state<=12;
					out<=148;
				end
				if(in == 718) begin
					state<=12;
					out<=149;
				end
				if(in == 719) begin
					state<=12;
					out<=150;
				end
				if(in == 720) begin
					state<=12;
					out<=151;
				end
				if(in == 721) begin
					state<=18;
					out<=152;
				end
				if(in == 722) begin
					state<=18;
					out<=153;
				end
				if(in == 723) begin
					state<=18;
					out<=154;
				end
				if(in == 724) begin
					state<=18;
					out<=155;
				end
				if(in == 725) begin
					state<=24;
					out<=156;
				end
				if(in == 726) begin
					state<=24;
					out<=157;
				end
				if(in == 727) begin
					state<=24;
					out<=158;
				end
				if(in == 728) begin
					state<=24;
					out<=159;
				end
				if(in == 729) begin
					state<=8;
					out<=160;
				end
				if(in == 730) begin
					state<=8;
					out<=161;
				end
				if(in == 731) begin
					state<=8;
					out<=162;
				end
				if(in == 732) begin
					state<=8;
					out<=163;
				end
				if(in == 733) begin
					state<=12;
					out<=164;
				end
				if(in == 734) begin
					state<=12;
					out<=165;
				end
				if(in == 735) begin
					state<=12;
					out<=166;
				end
				if(in == 736) begin
					state<=12;
					out<=167;
				end
				if(in == 737) begin
					state<=18;
					out<=168;
				end
				if(in == 738) begin
					state<=18;
					out<=169;
				end
				if(in == 739) begin
					state<=18;
					out<=170;
				end
				if(in == 740) begin
					state<=18;
					out<=171;
				end
				if(in == 741) begin
					state<=24;
					out<=172;
				end
				if(in == 742) begin
					state<=24;
					out<=173;
				end
				if(in == 743) begin
					state<=24;
					out<=174;
				end
				if(in == 744) begin
					state<=24;
					out<=175;
				end
				if(in == 745) begin
					state<=8;
					out<=176;
				end
				if(in == 746) begin
					state<=8;
					out<=177;
				end
				if(in == 747) begin
					state<=8;
					out<=178;
				end
				if(in == 748) begin
					state<=8;
					out<=179;
				end
				if(in == 749) begin
					state<=3;
					out<=180;
				end
				if(in == 750) begin
					state<=7;
					out<=181;
				end
				if(in == 751) begin
					state<=3;
					out<=182;
				end
				if(in == 752) begin
					state<=12;
					out<=183;
				end
				if(in == 753) begin
					state<=3;
					out<=184;
				end
				if(in == 754) begin
					state<=12;
					out<=185;
				end
				if(in == 755) begin
					state<=12;
					out<=186;
				end
				if(in == 756) begin
					state<=12;
					out<=187;
				end
				if(in == 757) begin
					state<=18;
					out<=188;
				end
				if(in == 758) begin
					state<=18;
					out<=189;
				end
				if(in == 759) begin
					state<=18;
					out<=190;
				end
				if(in == 760) begin
					state<=18;
					out<=191;
				end
				if(in == 761) begin
					state<=24;
					out<=192;
				end
				if(in == 762) begin
					state<=24;
					out<=193;
				end
				if(in == 763) begin
					state<=24;
					out<=194;
				end
				if(in == 764) begin
					state<=24;
					out<=195;
				end
				if(in == 765) begin
					state<=8;
					out<=196;
				end
				if(in == 766) begin
					state<=8;
					out<=197;
				end
				if(in == 767) begin
					state<=8;
					out<=198;
				end
				if(in == 768) begin
					state<=8;
					out<=199;
				end
				if(in == 769) begin
					state<=12;
					out<=200;
				end
				if(in == 770) begin
					state<=12;
					out<=201;
				end
				if(in == 771) begin
					state<=12;
					out<=202;
				end
				if(in == 772) begin
					state<=12;
					out<=203;
				end
				if(in == 773) begin
					state<=18;
					out<=204;
				end
				if(in == 774) begin
					state<=18;
					out<=205;
				end
				if(in == 775) begin
					state<=18;
					out<=206;
				end
				if(in == 776) begin
					state<=18;
					out<=207;
				end
				if(in == 777) begin
					state<=24;
					out<=208;
				end
				if(in == 778) begin
					state<=24;
					out<=209;
				end
				if(in == 779) begin
					state<=24;
					out<=210;
				end
				if(in == 780) begin
					state<=24;
					out<=211;
				end
				if(in == 781) begin
					state<=8;
					out<=212;
				end
				if(in == 782) begin
					state<=8;
					out<=213;
				end
				if(in == 783) begin
					state<=8;
					out<=214;
				end
				if(in == 784) begin
					state<=8;
					out<=215;
				end
				if(in == 785) begin
					state<=12;
					out<=216;
				end
				if(in == 786) begin
					state<=12;
					out<=217;
				end
				if(in == 787) begin
					state<=12;
					out<=218;
				end
				if(in == 788) begin
					state<=12;
					out<=219;
				end
				if(in == 789) begin
					state<=18;
					out<=220;
				end
				if(in == 790) begin
					state<=18;
					out<=221;
				end
				if(in == 791) begin
					state<=18;
					out<=222;
				end
				if(in == 792) begin
					state<=18;
					out<=223;
				end
				if(in == 793) begin
					state<=24;
					out<=224;
				end
				if(in == 794) begin
					state<=24;
					out<=225;
				end
				if(in == 795) begin
					state<=24;
					out<=226;
				end
				if(in == 796) begin
					state<=24;
					out<=227;
				end
				if(in == 797) begin
					state<=8;
					out<=228;
				end
				if(in == 798) begin
					state<=8;
					out<=229;
				end
				if(in == 799) begin
					state<=8;
					out<=230;
				end
				if(in == 800) begin
					state<=8;
					out<=231;
				end
				if(in == 801) begin
					state<=2;
					out<=232;
				end
				if(in == 802) begin
					state<=2;
					out<=233;
				end
				if(in == 803) begin
					state<=2;
					out<=234;
				end
				if(in == 804) begin
					state<=2;
					out<=235;
				end
				if(in == 805) begin
					state<=2;
					out<=236;
				end
				if(in == 806) begin
					state<=2;
					out<=237;
				end
				if(in == 807) begin
					state<=2;
					out<=238;
				end
				if(in == 808) begin
					state<=2;
					out<=239;
				end
				if(in == 809) begin
					state<=2;
					out<=240;
				end
				if(in == 810) begin
					state<=2;
					out<=241;
				end
				if(in == 811) begin
					state<=2;
					out<=242;
				end
				if(in == 812) begin
					state<=2;
					out<=243;
				end
				if(in == 813) begin
					state<=3;
					out<=244;
				end
				if(in == 814) begin
					state<=7;
					out<=245;
				end
				if(in == 815) begin
					state<=3;
					out<=246;
				end
				if(in == 816) begin
					state<=12;
					out<=247;
				end
				if(in == 817) begin
					state<=3;
					out<=248;
				end
				if(in == 818) begin
					state<=12;
					out<=249;
				end
				if(in == 819) begin
					state<=12;
					out<=250;
				end
				if(in == 820) begin
					state<=12;
					out<=251;
				end
				if(in == 821) begin
					state<=18;
					out<=252;
				end
				if(in == 822) begin
					state<=18;
					out<=253;
				end
				if(in == 823) begin
					state<=18;
					out<=254;
				end
				if(in == 824) begin
					state<=18;
					out<=255;
				end
				if(in == 825) begin
					state<=24;
					out<=0;
				end
				if(in == 826) begin
					state<=24;
					out<=1;
				end
				if(in == 827) begin
					state<=24;
					out<=2;
				end
				if(in == 828) begin
					state<=24;
					out<=3;
				end
				if(in == 829) begin
					state<=8;
					out<=4;
				end
				if(in == 830) begin
					state<=8;
					out<=5;
				end
				if(in == 831) begin
					state<=8;
					out<=6;
				end
				if(in == 832) begin
					state<=8;
					out<=7;
				end
				if(in == 833) begin
					state<=12;
					out<=8;
				end
				if(in == 834) begin
					state<=12;
					out<=9;
				end
				if(in == 835) begin
					state<=12;
					out<=10;
				end
				if(in == 836) begin
					state<=12;
					out<=11;
				end
				if(in == 837) begin
					state<=18;
					out<=12;
				end
				if(in == 838) begin
					state<=18;
					out<=13;
				end
				if(in == 839) begin
					state<=18;
					out<=14;
				end
				if(in == 840) begin
					state<=18;
					out<=15;
				end
				if(in == 841) begin
					state<=24;
					out<=16;
				end
				if(in == 842) begin
					state<=24;
					out<=17;
				end
				if(in == 843) begin
					state<=24;
					out<=18;
				end
				if(in == 844) begin
					state<=24;
					out<=19;
				end
				if(in == 845) begin
					state<=8;
					out<=20;
				end
				if(in == 846) begin
					state<=8;
					out<=21;
				end
				if(in == 847) begin
					state<=8;
					out<=22;
				end
				if(in == 848) begin
					state<=8;
					out<=23;
				end
				if(in == 849) begin
					state<=12;
					out<=24;
				end
				if(in == 850) begin
					state<=12;
					out<=25;
				end
				if(in == 851) begin
					state<=12;
					out<=26;
				end
				if(in == 852) begin
					state<=12;
					out<=27;
				end
				if(in == 853) begin
					state<=18;
					out<=28;
				end
				if(in == 854) begin
					state<=18;
					out<=29;
				end
				if(in == 855) begin
					state<=18;
					out<=30;
				end
				if(in == 856) begin
					state<=18;
					out<=31;
				end
				if(in == 857) begin
					state<=24;
					out<=32;
				end
				if(in == 858) begin
					state<=24;
					out<=33;
				end
				if(in == 859) begin
					state<=24;
					out<=34;
				end
				if(in == 860) begin
					state<=24;
					out<=35;
				end
				if(in == 861) begin
					state<=8;
					out<=36;
				end
				if(in == 862) begin
					state<=8;
					out<=37;
				end
				if(in == 863) begin
					state<=8;
					out<=38;
				end
				if(in == 864) begin
					state<=8;
					out<=39;
				end
				if(in == 865) begin
					state<=3;
					out<=40;
				end
				if(in == 866) begin
					state<=7;
					out<=41;
				end
				if(in == 867) begin
					state<=3;
					out<=42;
				end
				if(in == 868) begin
					state<=12;
					out<=43;
				end
				if(in == 869) begin
					state<=3;
					out<=44;
				end
				if(in == 870) begin
					state<=12;
					out<=45;
				end
				if(in == 871) begin
					state<=12;
					out<=46;
				end
				if(in == 872) begin
					state<=12;
					out<=47;
				end
				if(in == 873) begin
					state<=18;
					out<=48;
				end
				if(in == 874) begin
					state<=18;
					out<=49;
				end
				if(in == 875) begin
					state<=18;
					out<=50;
				end
				if(in == 876) begin
					state<=18;
					out<=51;
				end
				if(in == 877) begin
					state<=24;
					out<=52;
				end
				if(in == 878) begin
					state<=24;
					out<=53;
				end
				if(in == 879) begin
					state<=24;
					out<=54;
				end
				if(in == 880) begin
					state<=24;
					out<=55;
				end
				if(in == 881) begin
					state<=8;
					out<=56;
				end
				if(in == 882) begin
					state<=8;
					out<=57;
				end
				if(in == 883) begin
					state<=8;
					out<=58;
				end
				if(in == 884) begin
					state<=8;
					out<=59;
				end
				if(in == 885) begin
					state<=12;
					out<=60;
				end
				if(in == 886) begin
					state<=12;
					out<=61;
				end
				if(in == 887) begin
					state<=12;
					out<=62;
				end
				if(in == 888) begin
					state<=12;
					out<=63;
				end
				if(in == 889) begin
					state<=18;
					out<=64;
				end
				if(in == 890) begin
					state<=18;
					out<=65;
				end
				if(in == 891) begin
					state<=18;
					out<=66;
				end
				if(in == 892) begin
					state<=18;
					out<=67;
				end
				if(in == 893) begin
					state<=24;
					out<=68;
				end
				if(in == 894) begin
					state<=24;
					out<=69;
				end
				if(in == 895) begin
					state<=24;
					out<=70;
				end
				if(in == 896) begin
					state<=24;
					out<=71;
				end
				if(in == 897) begin
					state<=8;
					out<=72;
				end
				if(in == 898) begin
					state<=8;
					out<=73;
				end
				if(in == 899) begin
					state<=8;
					out<=74;
				end
				if(in == 900) begin
					state<=8;
					out<=75;
				end
				if(in == 901) begin
					state<=12;
					out<=76;
				end
				if(in == 902) begin
					state<=12;
					out<=77;
				end
				if(in == 903) begin
					state<=12;
					out<=78;
				end
				if(in == 904) begin
					state<=12;
					out<=79;
				end
				if(in == 905) begin
					state<=18;
					out<=80;
				end
				if(in == 906) begin
					state<=18;
					out<=81;
				end
				if(in == 907) begin
					state<=18;
					out<=82;
				end
				if(in == 908) begin
					state<=18;
					out<=83;
				end
				if(in == 909) begin
					state<=24;
					out<=84;
				end
				if(in == 910) begin
					state<=24;
					out<=85;
				end
				if(in == 911) begin
					state<=24;
					out<=86;
				end
				if(in == 912) begin
					state<=24;
					out<=87;
				end
				if(in == 913) begin
					state<=8;
					out<=88;
				end
				if(in == 914) begin
					state<=8;
					out<=89;
				end
				if(in == 915) begin
					state<=8;
					out<=90;
				end
				if(in == 916) begin
					state<=8;
					out<=91;
				end
				if(in == 917) begin
					state<=2;
					out<=92;
				end
				if(in == 918) begin
					state<=2;
					out<=93;
				end
				if(in == 919) begin
					state<=2;
					out<=94;
				end
				if(in == 920) begin
					state<=2;
					out<=95;
				end
				if(in == 921) begin
					state<=2;
					out<=96;
				end
				if(in == 922) begin
					state<=2;
					out<=97;
				end
				if(in == 923) begin
					state<=2;
					out<=98;
				end
				if(in == 924) begin
					state<=2;
					out<=99;
				end
				if(in == 925) begin
					state<=2;
					out<=100;
				end
				if(in == 926) begin
					state<=2;
					out<=101;
				end
				if(in == 927) begin
					state<=2;
					out<=102;
				end
				if(in == 928) begin
					state<=2;
					out<=103;
				end
			end
			8: begin
				if(in == 0) begin
					state<=3;
					out<=104;
				end
				if(in == 1) begin
					state<=1;
					out<=105;
				end
				if(in == 2) begin
					state<=8;
					out<=106;
				end
				if(in == 3) begin
					state<=3;
					out<=107;
				end
				if(in == 4) begin
					state<=12;
					out<=108;
				end
				if(in == 5) begin
					state<=3;
					out<=109;
				end
				if(in == 6) begin
					state<=12;
					out<=110;
				end
				if(in == 7) begin
					state<=9;
					out<=111;
				end
				if(in == 8) begin
					state<=9;
					out<=112;
				end
				if(in == 9) begin
					state<=12;
					out<=113;
				end
				if(in == 10) begin
					state<=12;
					out<=114;
				end
				if(in == 11) begin
					state<=9;
					out<=115;
				end
				if(in == 12) begin
					state<=9;
					out<=116;
				end
				if(in == 13) begin
					state<=12;
					out<=117;
				end
				if(in == 14) begin
					state<=12;
					out<=118;
				end
				if(in == 15) begin
					state<=9;
					out<=119;
				end
				if(in == 16) begin
					state<=9;
					out<=120;
				end
				if(in == 17) begin
					state<=12;
					out<=121;
				end
				if(in == 18) begin
					state<=12;
					out<=122;
				end
				if(in == 19) begin
					state<=9;
					out<=123;
				end
				if(in == 20) begin
					state<=9;
					out<=124;
				end
				if(in == 21) begin
					state<=12;
					out<=125;
				end
				if(in == 22) begin
					state<=12;
					out<=126;
				end
				if(in == 23) begin
					state<=9;
					out<=127;
				end
				if(in == 24) begin
					state<=9;
					out<=128;
				end
				if(in == 25) begin
					state<=12;
					out<=129;
				end
				if(in == 26) begin
					state<=12;
					out<=130;
				end
				if(in == 27) begin
					state<=9;
					out<=131;
				end
				if(in == 28) begin
					state<=9;
					out<=132;
				end
				if(in == 29) begin
					state<=12;
					out<=133;
				end
				if(in == 30) begin
					state<=12;
					out<=134;
				end
				if(in == 31) begin
					state<=9;
					out<=135;
				end
				if(in == 32) begin
					state<=9;
					out<=136;
				end
				if(in == 33) begin
					state<=12;
					out<=137;
				end
				if(in == 34) begin
					state<=12;
					out<=138;
				end
				if(in == 35) begin
					state<=9;
					out<=139;
				end
				if(in == 36) begin
					state<=9;
					out<=140;
				end
				if(in == 37) begin
					state<=12;
					out<=141;
				end
				if(in == 38) begin
					state<=12;
					out<=142;
				end
				if(in == 39) begin
					state<=9;
					out<=143;
				end
				if(in == 40) begin
					state<=9;
					out<=144;
				end
				if(in == 41) begin
					state<=12;
					out<=145;
				end
				if(in == 42) begin
					state<=12;
					out<=146;
				end
				if(in == 43) begin
					state<=9;
					out<=147;
				end
				if(in == 44) begin
					state<=9;
					out<=148;
				end
				if(in == 45) begin
					state<=12;
					out<=149;
				end
				if(in == 46) begin
					state<=12;
					out<=150;
				end
				if(in == 47) begin
					state<=9;
					out<=151;
				end
				if(in == 48) begin
					state<=9;
					out<=152;
				end
				if(in == 49) begin
					state<=12;
					out<=153;
				end
				if(in == 50) begin
					state<=12;
					out<=154;
				end
				if(in == 51) begin
					state<=9;
					out<=155;
				end
				if(in == 52) begin
					state<=9;
					out<=156;
				end
				if(in == 53) begin
					state<=3;
					out<=157;
				end
				if(in == 54) begin
					state<=8;
					out<=158;
				end
				if(in == 55) begin
					state<=3;
					out<=159;
				end
				if(in == 56) begin
					state<=12;
					out<=160;
				end
				if(in == 57) begin
					state<=3;
					out<=161;
				end
				if(in == 58) begin
					state<=12;
					out<=162;
				end
				if(in == 59) begin
					state<=9;
					out<=163;
				end
				if(in == 60) begin
					state<=9;
					out<=164;
				end
				if(in == 61) begin
					state<=12;
					out<=165;
				end
				if(in == 62) begin
					state<=12;
					out<=166;
				end
				if(in == 63) begin
					state<=9;
					out<=167;
				end
				if(in == 64) begin
					state<=9;
					out<=168;
				end
				if(in == 65) begin
					state<=12;
					out<=169;
				end
				if(in == 66) begin
					state<=12;
					out<=170;
				end
				if(in == 67) begin
					state<=9;
					out<=171;
				end
				if(in == 68) begin
					state<=9;
					out<=172;
				end
				if(in == 69) begin
					state<=12;
					out<=173;
				end
				if(in == 70) begin
					state<=12;
					out<=174;
				end
				if(in == 71) begin
					state<=9;
					out<=175;
				end
				if(in == 72) begin
					state<=9;
					out<=176;
				end
				if(in == 73) begin
					state<=12;
					out<=177;
				end
				if(in == 74) begin
					state<=12;
					out<=178;
				end
				if(in == 75) begin
					state<=9;
					out<=179;
				end
				if(in == 76) begin
					state<=9;
					out<=180;
				end
				if(in == 77) begin
					state<=12;
					out<=181;
				end
				if(in == 78) begin
					state<=12;
					out<=182;
				end
				if(in == 79) begin
					state<=9;
					out<=183;
				end
				if(in == 80) begin
					state<=9;
					out<=184;
				end
				if(in == 81) begin
					state<=12;
					out<=185;
				end
				if(in == 82) begin
					state<=12;
					out<=186;
				end
				if(in == 83) begin
					state<=9;
					out<=187;
				end
				if(in == 84) begin
					state<=9;
					out<=188;
				end
				if(in == 85) begin
					state<=12;
					out<=189;
				end
				if(in == 86) begin
					state<=12;
					out<=190;
				end
				if(in == 87) begin
					state<=9;
					out<=191;
				end
				if(in == 88) begin
					state<=9;
					out<=192;
				end
				if(in == 89) begin
					state<=12;
					out<=193;
				end
				if(in == 90) begin
					state<=12;
					out<=194;
				end
				if(in == 91) begin
					state<=9;
					out<=195;
				end
				if(in == 92) begin
					state<=9;
					out<=196;
				end
				if(in == 93) begin
					state<=12;
					out<=197;
				end
				if(in == 94) begin
					state<=12;
					out<=198;
				end
				if(in == 95) begin
					state<=9;
					out<=199;
				end
				if(in == 96) begin
					state<=9;
					out<=200;
				end
				if(in == 97) begin
					state<=12;
					out<=201;
				end
				if(in == 98) begin
					state<=12;
					out<=202;
				end
				if(in == 99) begin
					state<=9;
					out<=203;
				end
				if(in == 100) begin
					state<=9;
					out<=204;
				end
				if(in == 101) begin
					state<=12;
					out<=205;
				end
				if(in == 102) begin
					state<=12;
					out<=206;
				end
				if(in == 103) begin
					state<=9;
					out<=207;
				end
				if(in == 104) begin
					state<=9;
					out<=208;
				end
				if(in == 105) begin
					state<=2;
					out<=209;
				end
				if(in == 106) begin
					state<=2;
					out<=210;
				end
				if(in == 107) begin
					state<=2;
					out<=211;
				end
				if(in == 108) begin
					state<=2;
					out<=212;
				end
				if(in == 109) begin
					state<=2;
					out<=213;
				end
				if(in == 110) begin
					state<=2;
					out<=214;
				end
				if(in == 111) begin
					state<=2;
					out<=215;
				end
				if(in == 112) begin
					state<=2;
					out<=216;
				end
				if(in == 113) begin
					state<=2;
					out<=217;
				end
				if(in == 114) begin
					state<=2;
					out<=218;
				end
				if(in == 115) begin
					state<=2;
					out<=219;
				end
				if(in == 116) begin
					state<=2;
					out<=220;
				end
				if(in == 117) begin
					state<=3;
					out<=221;
				end
				if(in == 118) begin
					state<=8;
					out<=222;
				end
				if(in == 119) begin
					state<=3;
					out<=223;
				end
				if(in == 120) begin
					state<=12;
					out<=224;
				end
				if(in == 121) begin
					state<=3;
					out<=225;
				end
				if(in == 122) begin
					state<=12;
					out<=226;
				end
				if(in == 123) begin
					state<=9;
					out<=227;
				end
				if(in == 124) begin
					state<=9;
					out<=228;
				end
				if(in == 125) begin
					state<=12;
					out<=229;
				end
				if(in == 126) begin
					state<=12;
					out<=230;
				end
				if(in == 127) begin
					state<=9;
					out<=231;
				end
				if(in == 128) begin
					state<=9;
					out<=232;
				end
				if(in == 129) begin
					state<=12;
					out<=233;
				end
				if(in == 130) begin
					state<=12;
					out<=234;
				end
				if(in == 131) begin
					state<=9;
					out<=235;
				end
				if(in == 132) begin
					state<=9;
					out<=236;
				end
				if(in == 133) begin
					state<=12;
					out<=237;
				end
				if(in == 134) begin
					state<=12;
					out<=238;
				end
				if(in == 135) begin
					state<=9;
					out<=239;
				end
				if(in == 136) begin
					state<=9;
					out<=240;
				end
				if(in == 137) begin
					state<=12;
					out<=241;
				end
				if(in == 138) begin
					state<=12;
					out<=242;
				end
				if(in == 139) begin
					state<=9;
					out<=243;
				end
				if(in == 140) begin
					state<=9;
					out<=244;
				end
				if(in == 141) begin
					state<=12;
					out<=245;
				end
				if(in == 142) begin
					state<=12;
					out<=246;
				end
				if(in == 143) begin
					state<=9;
					out<=247;
				end
				if(in == 144) begin
					state<=9;
					out<=248;
				end
				if(in == 145) begin
					state<=12;
					out<=249;
				end
				if(in == 146) begin
					state<=12;
					out<=250;
				end
				if(in == 147) begin
					state<=9;
					out<=251;
				end
				if(in == 148) begin
					state<=9;
					out<=252;
				end
				if(in == 149) begin
					state<=12;
					out<=253;
				end
				if(in == 150) begin
					state<=12;
					out<=254;
				end
				if(in == 151) begin
					state<=9;
					out<=255;
				end
				if(in == 152) begin
					state<=9;
					out<=0;
				end
				if(in == 153) begin
					state<=12;
					out<=1;
				end
				if(in == 154) begin
					state<=12;
					out<=2;
				end
				if(in == 155) begin
					state<=9;
					out<=3;
				end
				if(in == 156) begin
					state<=9;
					out<=4;
				end
				if(in == 157) begin
					state<=12;
					out<=5;
				end
				if(in == 158) begin
					state<=12;
					out<=6;
				end
				if(in == 159) begin
					state<=9;
					out<=7;
				end
				if(in == 160) begin
					state<=9;
					out<=8;
				end
				if(in == 161) begin
					state<=12;
					out<=9;
				end
				if(in == 162) begin
					state<=12;
					out<=10;
				end
				if(in == 163) begin
					state<=9;
					out<=11;
				end
				if(in == 164) begin
					state<=9;
					out<=12;
				end
				if(in == 165) begin
					state<=12;
					out<=13;
				end
				if(in == 166) begin
					state<=12;
					out<=14;
				end
				if(in == 167) begin
					state<=9;
					out<=15;
				end
				if(in == 168) begin
					state<=9;
					out<=16;
				end
				if(in == 169) begin
					state<=3;
					out<=17;
				end
				if(in == 170) begin
					state<=8;
					out<=18;
				end
				if(in == 171) begin
					state<=3;
					out<=19;
				end
				if(in == 172) begin
					state<=12;
					out<=20;
				end
				if(in == 173) begin
					state<=3;
					out<=21;
				end
				if(in == 174) begin
					state<=12;
					out<=22;
				end
				if(in == 175) begin
					state<=9;
					out<=23;
				end
				if(in == 176) begin
					state<=9;
					out<=24;
				end
				if(in == 177) begin
					state<=12;
					out<=25;
				end
				if(in == 178) begin
					state<=12;
					out<=26;
				end
				if(in == 179) begin
					state<=9;
					out<=27;
				end
				if(in == 180) begin
					state<=9;
					out<=28;
				end
				if(in == 181) begin
					state<=12;
					out<=29;
				end
				if(in == 182) begin
					state<=12;
					out<=30;
				end
				if(in == 183) begin
					state<=9;
					out<=31;
				end
				if(in == 184) begin
					state<=9;
					out<=32;
				end
				if(in == 185) begin
					state<=12;
					out<=33;
				end
				if(in == 186) begin
					state<=12;
					out<=34;
				end
				if(in == 187) begin
					state<=9;
					out<=35;
				end
				if(in == 188) begin
					state<=9;
					out<=36;
				end
				if(in == 189) begin
					state<=12;
					out<=37;
				end
				if(in == 190) begin
					state<=12;
					out<=38;
				end
				if(in == 191) begin
					state<=9;
					out<=39;
				end
				if(in == 192) begin
					state<=9;
					out<=40;
				end
				if(in == 193) begin
					state<=12;
					out<=41;
				end
				if(in == 194) begin
					state<=12;
					out<=42;
				end
				if(in == 195) begin
					state<=9;
					out<=43;
				end
				if(in == 196) begin
					state<=9;
					out<=44;
				end
				if(in == 197) begin
					state<=12;
					out<=45;
				end
				if(in == 198) begin
					state<=12;
					out<=46;
				end
				if(in == 199) begin
					state<=9;
					out<=47;
				end
				if(in == 200) begin
					state<=9;
					out<=48;
				end
				if(in == 201) begin
					state<=12;
					out<=49;
				end
				if(in == 202) begin
					state<=12;
					out<=50;
				end
				if(in == 203) begin
					state<=9;
					out<=51;
				end
				if(in == 204) begin
					state<=9;
					out<=52;
				end
				if(in == 205) begin
					state<=12;
					out<=53;
				end
				if(in == 206) begin
					state<=12;
					out<=54;
				end
				if(in == 207) begin
					state<=9;
					out<=55;
				end
				if(in == 208) begin
					state<=9;
					out<=56;
				end
				if(in == 209) begin
					state<=12;
					out<=57;
				end
				if(in == 210) begin
					state<=12;
					out<=58;
				end
				if(in == 211) begin
					state<=9;
					out<=59;
				end
				if(in == 212) begin
					state<=9;
					out<=60;
				end
				if(in == 213) begin
					state<=12;
					out<=61;
				end
				if(in == 214) begin
					state<=12;
					out<=62;
				end
				if(in == 215) begin
					state<=9;
					out<=63;
				end
				if(in == 216) begin
					state<=9;
					out<=64;
				end
				if(in == 217) begin
					state<=12;
					out<=65;
				end
				if(in == 218) begin
					state<=12;
					out<=66;
				end
				if(in == 219) begin
					state<=9;
					out<=67;
				end
				if(in == 220) begin
					state<=9;
					out<=68;
				end
				if(in == 221) begin
					state<=2;
					out<=69;
				end
				if(in == 222) begin
					state<=2;
					out<=70;
				end
				if(in == 223) begin
					state<=2;
					out<=71;
				end
				if(in == 224) begin
					state<=2;
					out<=72;
				end
				if(in == 225) begin
					state<=2;
					out<=73;
				end
				if(in == 226) begin
					state<=2;
					out<=74;
				end
				if(in == 227) begin
					state<=2;
					out<=75;
				end
				if(in == 228) begin
					state<=2;
					out<=76;
				end
				if(in == 229) begin
					state<=2;
					out<=77;
				end
				if(in == 230) begin
					state<=2;
					out<=78;
				end
				if(in == 231) begin
					state<=2;
					out<=79;
				end
				if(in == 232) begin
					state<=2;
					out<=80;
				end
				if(in == 233) begin
					state<=3;
					out<=81;
				end
				if(in == 234) begin
					state<=8;
					out<=82;
				end
				if(in == 235) begin
					state<=3;
					out<=83;
				end
				if(in == 236) begin
					state<=12;
					out<=84;
				end
				if(in == 237) begin
					state<=3;
					out<=85;
				end
				if(in == 238) begin
					state<=12;
					out<=86;
				end
				if(in == 239) begin
					state<=9;
					out<=87;
				end
				if(in == 240) begin
					state<=9;
					out<=88;
				end
				if(in == 241) begin
					state<=12;
					out<=89;
				end
				if(in == 242) begin
					state<=12;
					out<=90;
				end
				if(in == 243) begin
					state<=9;
					out<=91;
				end
				if(in == 244) begin
					state<=9;
					out<=92;
				end
				if(in == 245) begin
					state<=12;
					out<=93;
				end
				if(in == 246) begin
					state<=12;
					out<=94;
				end
				if(in == 247) begin
					state<=9;
					out<=95;
				end
				if(in == 248) begin
					state<=9;
					out<=96;
				end
				if(in == 249) begin
					state<=12;
					out<=97;
				end
				if(in == 250) begin
					state<=12;
					out<=98;
				end
				if(in == 251) begin
					state<=9;
					out<=99;
				end
				if(in == 252) begin
					state<=9;
					out<=100;
				end
				if(in == 253) begin
					state<=12;
					out<=101;
				end
				if(in == 254) begin
					state<=12;
					out<=102;
				end
				if(in == 255) begin
					state<=9;
					out<=103;
				end
				if(in == 256) begin
					state<=9;
					out<=104;
				end
				if(in == 257) begin
					state<=12;
					out<=105;
				end
				if(in == 258) begin
					state<=12;
					out<=106;
				end
				if(in == 259) begin
					state<=9;
					out<=107;
				end
				if(in == 260) begin
					state<=9;
					out<=108;
				end
				if(in == 261) begin
					state<=12;
					out<=109;
				end
				if(in == 262) begin
					state<=12;
					out<=110;
				end
				if(in == 263) begin
					state<=9;
					out<=111;
				end
				if(in == 264) begin
					state<=9;
					out<=112;
				end
				if(in == 265) begin
					state<=12;
					out<=113;
				end
				if(in == 266) begin
					state<=12;
					out<=114;
				end
				if(in == 267) begin
					state<=9;
					out<=115;
				end
				if(in == 268) begin
					state<=9;
					out<=116;
				end
				if(in == 269) begin
					state<=12;
					out<=117;
				end
				if(in == 270) begin
					state<=12;
					out<=118;
				end
				if(in == 271) begin
					state<=9;
					out<=119;
				end
				if(in == 272) begin
					state<=9;
					out<=120;
				end
				if(in == 273) begin
					state<=12;
					out<=121;
				end
				if(in == 274) begin
					state<=12;
					out<=122;
				end
				if(in == 275) begin
					state<=9;
					out<=123;
				end
				if(in == 276) begin
					state<=9;
					out<=124;
				end
				if(in == 277) begin
					state<=12;
					out<=125;
				end
				if(in == 278) begin
					state<=12;
					out<=126;
				end
				if(in == 279) begin
					state<=9;
					out<=127;
				end
				if(in == 280) begin
					state<=9;
					out<=128;
				end
				if(in == 281) begin
					state<=12;
					out<=129;
				end
				if(in == 282) begin
					state<=12;
					out<=130;
				end
				if(in == 283) begin
					state<=9;
					out<=131;
				end
				if(in == 284) begin
					state<=9;
					out<=132;
				end
				if(in == 285) begin
					state<=3;
					out<=133;
				end
				if(in == 286) begin
					state<=8;
					out<=134;
				end
				if(in == 287) begin
					state<=3;
					out<=135;
				end
				if(in == 288) begin
					state<=12;
					out<=136;
				end
				if(in == 289) begin
					state<=3;
					out<=137;
				end
				if(in == 290) begin
					state<=12;
					out<=138;
				end
				if(in == 291) begin
					state<=9;
					out<=139;
				end
				if(in == 292) begin
					state<=9;
					out<=140;
				end
				if(in == 293) begin
					state<=12;
					out<=141;
				end
				if(in == 294) begin
					state<=12;
					out<=142;
				end
				if(in == 295) begin
					state<=9;
					out<=143;
				end
				if(in == 296) begin
					state<=9;
					out<=144;
				end
				if(in == 297) begin
					state<=12;
					out<=145;
				end
				if(in == 298) begin
					state<=12;
					out<=146;
				end
				if(in == 299) begin
					state<=9;
					out<=147;
				end
				if(in == 300) begin
					state<=9;
					out<=148;
				end
				if(in == 301) begin
					state<=12;
					out<=149;
				end
				if(in == 302) begin
					state<=12;
					out<=150;
				end
				if(in == 303) begin
					state<=9;
					out<=151;
				end
				if(in == 304) begin
					state<=9;
					out<=152;
				end
				if(in == 305) begin
					state<=12;
					out<=153;
				end
				if(in == 306) begin
					state<=12;
					out<=154;
				end
				if(in == 307) begin
					state<=9;
					out<=155;
				end
				if(in == 308) begin
					state<=9;
					out<=156;
				end
				if(in == 309) begin
					state<=12;
					out<=157;
				end
				if(in == 310) begin
					state<=12;
					out<=158;
				end
				if(in == 311) begin
					state<=9;
					out<=159;
				end
				if(in == 312) begin
					state<=9;
					out<=160;
				end
				if(in == 313) begin
					state<=12;
					out<=161;
				end
				if(in == 314) begin
					state<=12;
					out<=162;
				end
				if(in == 315) begin
					state<=9;
					out<=163;
				end
				if(in == 316) begin
					state<=9;
					out<=164;
				end
				if(in == 317) begin
					state<=12;
					out<=165;
				end
				if(in == 318) begin
					state<=12;
					out<=166;
				end
				if(in == 319) begin
					state<=9;
					out<=167;
				end
				if(in == 320) begin
					state<=9;
					out<=168;
				end
				if(in == 321) begin
					state<=12;
					out<=169;
				end
				if(in == 322) begin
					state<=12;
					out<=170;
				end
				if(in == 323) begin
					state<=9;
					out<=171;
				end
				if(in == 324) begin
					state<=9;
					out<=172;
				end
				if(in == 325) begin
					state<=12;
					out<=173;
				end
				if(in == 326) begin
					state<=12;
					out<=174;
				end
				if(in == 327) begin
					state<=9;
					out<=175;
				end
				if(in == 328) begin
					state<=9;
					out<=176;
				end
				if(in == 329) begin
					state<=12;
					out<=177;
				end
				if(in == 330) begin
					state<=12;
					out<=178;
				end
				if(in == 331) begin
					state<=9;
					out<=179;
				end
				if(in == 332) begin
					state<=9;
					out<=180;
				end
				if(in == 333) begin
					state<=12;
					out<=181;
				end
				if(in == 334) begin
					state<=12;
					out<=182;
				end
				if(in == 335) begin
					state<=9;
					out<=183;
				end
				if(in == 336) begin
					state<=9;
					out<=184;
				end
				if(in == 337) begin
					state<=2;
					out<=185;
				end
				if(in == 338) begin
					state<=2;
					out<=186;
				end
				if(in == 339) begin
					state<=2;
					out<=187;
				end
				if(in == 340) begin
					state<=2;
					out<=188;
				end
				if(in == 341) begin
					state<=2;
					out<=189;
				end
				if(in == 342) begin
					state<=2;
					out<=190;
				end
				if(in == 343) begin
					state<=2;
					out<=191;
				end
				if(in == 344) begin
					state<=2;
					out<=192;
				end
				if(in == 345) begin
					state<=2;
					out<=193;
				end
				if(in == 346) begin
					state<=2;
					out<=194;
				end
				if(in == 347) begin
					state<=2;
					out<=195;
				end
				if(in == 348) begin
					state<=2;
					out<=196;
				end
				if(in == 349) begin
					state<=3;
					out<=197;
				end
				if(in == 350) begin
					state<=8;
					out<=198;
				end
				if(in == 351) begin
					state<=3;
					out<=199;
				end
				if(in == 352) begin
					state<=12;
					out<=200;
				end
				if(in == 353) begin
					state<=3;
					out<=201;
				end
				if(in == 354) begin
					state<=12;
					out<=202;
				end
				if(in == 355) begin
					state<=9;
					out<=203;
				end
				if(in == 356) begin
					state<=9;
					out<=204;
				end
				if(in == 357) begin
					state<=12;
					out<=205;
				end
				if(in == 358) begin
					state<=12;
					out<=206;
				end
				if(in == 359) begin
					state<=9;
					out<=207;
				end
				if(in == 360) begin
					state<=9;
					out<=208;
				end
				if(in == 361) begin
					state<=12;
					out<=209;
				end
				if(in == 362) begin
					state<=12;
					out<=210;
				end
				if(in == 363) begin
					state<=9;
					out<=211;
				end
				if(in == 364) begin
					state<=9;
					out<=212;
				end
				if(in == 365) begin
					state<=12;
					out<=213;
				end
				if(in == 366) begin
					state<=12;
					out<=214;
				end
				if(in == 367) begin
					state<=9;
					out<=215;
				end
				if(in == 368) begin
					state<=9;
					out<=216;
				end
				if(in == 369) begin
					state<=12;
					out<=217;
				end
				if(in == 370) begin
					state<=12;
					out<=218;
				end
				if(in == 371) begin
					state<=9;
					out<=219;
				end
				if(in == 372) begin
					state<=9;
					out<=220;
				end
				if(in == 373) begin
					state<=12;
					out<=221;
				end
				if(in == 374) begin
					state<=12;
					out<=222;
				end
				if(in == 375) begin
					state<=9;
					out<=223;
				end
				if(in == 376) begin
					state<=9;
					out<=224;
				end
				if(in == 377) begin
					state<=12;
					out<=225;
				end
				if(in == 378) begin
					state<=12;
					out<=226;
				end
				if(in == 379) begin
					state<=9;
					out<=227;
				end
				if(in == 380) begin
					state<=9;
					out<=228;
				end
				if(in == 381) begin
					state<=12;
					out<=229;
				end
				if(in == 382) begin
					state<=12;
					out<=230;
				end
				if(in == 383) begin
					state<=9;
					out<=231;
				end
				if(in == 384) begin
					state<=9;
					out<=232;
				end
				if(in == 385) begin
					state<=12;
					out<=233;
				end
				if(in == 386) begin
					state<=12;
					out<=234;
				end
				if(in == 387) begin
					state<=9;
					out<=235;
				end
				if(in == 388) begin
					state<=9;
					out<=236;
				end
				if(in == 389) begin
					state<=12;
					out<=237;
				end
				if(in == 390) begin
					state<=12;
					out<=238;
				end
				if(in == 391) begin
					state<=9;
					out<=239;
				end
				if(in == 392) begin
					state<=9;
					out<=240;
				end
				if(in == 393) begin
					state<=12;
					out<=241;
				end
				if(in == 394) begin
					state<=12;
					out<=242;
				end
				if(in == 395) begin
					state<=9;
					out<=243;
				end
				if(in == 396) begin
					state<=9;
					out<=244;
				end
				if(in == 397) begin
					state<=12;
					out<=245;
				end
				if(in == 398) begin
					state<=12;
					out<=246;
				end
				if(in == 399) begin
					state<=9;
					out<=247;
				end
				if(in == 400) begin
					state<=9;
					out<=248;
				end
				if(in == 401) begin
					state<=3;
					out<=249;
				end
				if(in == 402) begin
					state<=8;
					out<=250;
				end
				if(in == 403) begin
					state<=3;
					out<=251;
				end
				if(in == 404) begin
					state<=12;
					out<=252;
				end
				if(in == 405) begin
					state<=3;
					out<=253;
				end
				if(in == 406) begin
					state<=12;
					out<=254;
				end
				if(in == 407) begin
					state<=9;
					out<=255;
				end
				if(in == 408) begin
					state<=9;
					out<=0;
				end
				if(in == 409) begin
					state<=12;
					out<=1;
				end
				if(in == 410) begin
					state<=12;
					out<=2;
				end
				if(in == 411) begin
					state<=9;
					out<=3;
				end
				if(in == 412) begin
					state<=9;
					out<=4;
				end
				if(in == 413) begin
					state<=12;
					out<=5;
				end
				if(in == 414) begin
					state<=12;
					out<=6;
				end
				if(in == 415) begin
					state<=9;
					out<=7;
				end
				if(in == 416) begin
					state<=9;
					out<=8;
				end
				if(in == 417) begin
					state<=12;
					out<=9;
				end
				if(in == 418) begin
					state<=12;
					out<=10;
				end
				if(in == 419) begin
					state<=9;
					out<=11;
				end
				if(in == 420) begin
					state<=9;
					out<=12;
				end
				if(in == 421) begin
					state<=12;
					out<=13;
				end
				if(in == 422) begin
					state<=12;
					out<=14;
				end
				if(in == 423) begin
					state<=9;
					out<=15;
				end
				if(in == 424) begin
					state<=9;
					out<=16;
				end
				if(in == 425) begin
					state<=12;
					out<=17;
				end
				if(in == 426) begin
					state<=12;
					out<=18;
				end
				if(in == 427) begin
					state<=9;
					out<=19;
				end
				if(in == 428) begin
					state<=9;
					out<=20;
				end
				if(in == 429) begin
					state<=12;
					out<=21;
				end
				if(in == 430) begin
					state<=12;
					out<=22;
				end
				if(in == 431) begin
					state<=9;
					out<=23;
				end
				if(in == 432) begin
					state<=9;
					out<=24;
				end
				if(in == 433) begin
					state<=12;
					out<=25;
				end
				if(in == 434) begin
					state<=12;
					out<=26;
				end
				if(in == 435) begin
					state<=9;
					out<=27;
				end
				if(in == 436) begin
					state<=9;
					out<=28;
				end
				if(in == 437) begin
					state<=12;
					out<=29;
				end
				if(in == 438) begin
					state<=12;
					out<=30;
				end
				if(in == 439) begin
					state<=9;
					out<=31;
				end
				if(in == 440) begin
					state<=9;
					out<=32;
				end
				if(in == 441) begin
					state<=12;
					out<=33;
				end
				if(in == 442) begin
					state<=12;
					out<=34;
				end
				if(in == 443) begin
					state<=9;
					out<=35;
				end
				if(in == 444) begin
					state<=9;
					out<=36;
				end
				if(in == 445) begin
					state<=12;
					out<=37;
				end
				if(in == 446) begin
					state<=12;
					out<=38;
				end
				if(in == 447) begin
					state<=9;
					out<=39;
				end
				if(in == 448) begin
					state<=9;
					out<=40;
				end
				if(in == 449) begin
					state<=12;
					out<=41;
				end
				if(in == 450) begin
					state<=12;
					out<=42;
				end
				if(in == 451) begin
					state<=9;
					out<=43;
				end
				if(in == 452) begin
					state<=9;
					out<=44;
				end
				if(in == 453) begin
					state<=2;
					out<=45;
				end
				if(in == 454) begin
					state<=2;
					out<=46;
				end
				if(in == 455) begin
					state<=2;
					out<=47;
				end
				if(in == 456) begin
					state<=2;
					out<=48;
				end
				if(in == 457) begin
					state<=2;
					out<=49;
				end
				if(in == 458) begin
					state<=2;
					out<=50;
				end
				if(in == 459) begin
					state<=2;
					out<=51;
				end
				if(in == 460) begin
					state<=2;
					out<=52;
				end
				if(in == 461) begin
					state<=2;
					out<=53;
				end
				if(in == 462) begin
					state<=2;
					out<=54;
				end
				if(in == 463) begin
					state<=2;
					out<=55;
				end
				if(in == 464) begin
					state<=2;
					out<=56;
				end
				if(in == 465) begin
					state<=3;
					out<=57;
				end
				if(in == 466) begin
					state<=8;
					out<=58;
				end
				if(in == 467) begin
					state<=3;
					out<=59;
				end
				if(in == 468) begin
					state<=12;
					out<=60;
				end
				if(in == 469) begin
					state<=3;
					out<=61;
				end
				if(in == 470) begin
					state<=12;
					out<=62;
				end
				if(in == 471) begin
					state<=9;
					out<=63;
				end
				if(in == 472) begin
					state<=9;
					out<=64;
				end
				if(in == 473) begin
					state<=12;
					out<=65;
				end
				if(in == 474) begin
					state<=12;
					out<=66;
				end
				if(in == 475) begin
					state<=9;
					out<=67;
				end
				if(in == 476) begin
					state<=9;
					out<=68;
				end
				if(in == 477) begin
					state<=12;
					out<=69;
				end
				if(in == 478) begin
					state<=12;
					out<=70;
				end
				if(in == 479) begin
					state<=9;
					out<=71;
				end
				if(in == 480) begin
					state<=9;
					out<=72;
				end
				if(in == 481) begin
					state<=12;
					out<=73;
				end
				if(in == 482) begin
					state<=12;
					out<=74;
				end
				if(in == 483) begin
					state<=9;
					out<=75;
				end
				if(in == 484) begin
					state<=9;
					out<=76;
				end
				if(in == 485) begin
					state<=12;
					out<=77;
				end
				if(in == 486) begin
					state<=12;
					out<=78;
				end
				if(in == 487) begin
					state<=9;
					out<=79;
				end
				if(in == 488) begin
					state<=9;
					out<=80;
				end
				if(in == 489) begin
					state<=12;
					out<=81;
				end
				if(in == 490) begin
					state<=12;
					out<=82;
				end
				if(in == 491) begin
					state<=9;
					out<=83;
				end
				if(in == 492) begin
					state<=9;
					out<=84;
				end
				if(in == 493) begin
					state<=12;
					out<=85;
				end
				if(in == 494) begin
					state<=12;
					out<=86;
				end
				if(in == 495) begin
					state<=9;
					out<=87;
				end
				if(in == 496) begin
					state<=9;
					out<=88;
				end
				if(in == 497) begin
					state<=12;
					out<=89;
				end
				if(in == 498) begin
					state<=12;
					out<=90;
				end
				if(in == 499) begin
					state<=9;
					out<=91;
				end
				if(in == 500) begin
					state<=9;
					out<=92;
				end
				if(in == 501) begin
					state<=12;
					out<=93;
				end
				if(in == 502) begin
					state<=12;
					out<=94;
				end
				if(in == 503) begin
					state<=9;
					out<=95;
				end
				if(in == 504) begin
					state<=9;
					out<=96;
				end
				if(in == 505) begin
					state<=12;
					out<=97;
				end
				if(in == 506) begin
					state<=12;
					out<=98;
				end
				if(in == 507) begin
					state<=9;
					out<=99;
				end
				if(in == 508) begin
					state<=9;
					out<=100;
				end
				if(in == 509) begin
					state<=12;
					out<=101;
				end
				if(in == 510) begin
					state<=12;
					out<=102;
				end
				if(in == 511) begin
					state<=9;
					out<=103;
				end
				if(in == 512) begin
					state<=9;
					out<=104;
				end
				if(in == 513) begin
					state<=12;
					out<=105;
				end
				if(in == 514) begin
					state<=12;
					out<=106;
				end
				if(in == 515) begin
					state<=9;
					out<=107;
				end
				if(in == 516) begin
					state<=9;
					out<=108;
				end
				if(in == 517) begin
					state<=3;
					out<=109;
				end
				if(in == 518) begin
					state<=8;
					out<=110;
				end
				if(in == 519) begin
					state<=3;
					out<=111;
				end
				if(in == 520) begin
					state<=12;
					out<=112;
				end
				if(in == 521) begin
					state<=3;
					out<=113;
				end
				if(in == 522) begin
					state<=12;
					out<=114;
				end
				if(in == 523) begin
					state<=9;
					out<=115;
				end
				if(in == 524) begin
					state<=9;
					out<=116;
				end
				if(in == 525) begin
					state<=12;
					out<=117;
				end
				if(in == 526) begin
					state<=12;
					out<=118;
				end
				if(in == 527) begin
					state<=9;
					out<=119;
				end
				if(in == 528) begin
					state<=9;
					out<=120;
				end
				if(in == 529) begin
					state<=12;
					out<=121;
				end
				if(in == 530) begin
					state<=12;
					out<=122;
				end
				if(in == 531) begin
					state<=9;
					out<=123;
				end
				if(in == 532) begin
					state<=9;
					out<=124;
				end
				if(in == 533) begin
					state<=12;
					out<=125;
				end
				if(in == 534) begin
					state<=12;
					out<=126;
				end
				if(in == 535) begin
					state<=9;
					out<=127;
				end
				if(in == 536) begin
					state<=9;
					out<=128;
				end
				if(in == 537) begin
					state<=12;
					out<=129;
				end
				if(in == 538) begin
					state<=12;
					out<=130;
				end
				if(in == 539) begin
					state<=9;
					out<=131;
				end
				if(in == 540) begin
					state<=9;
					out<=132;
				end
				if(in == 541) begin
					state<=12;
					out<=133;
				end
				if(in == 542) begin
					state<=12;
					out<=134;
				end
				if(in == 543) begin
					state<=9;
					out<=135;
				end
				if(in == 544) begin
					state<=9;
					out<=136;
				end
				if(in == 545) begin
					state<=12;
					out<=137;
				end
				if(in == 546) begin
					state<=12;
					out<=138;
				end
				if(in == 547) begin
					state<=9;
					out<=139;
				end
				if(in == 548) begin
					state<=9;
					out<=140;
				end
				if(in == 549) begin
					state<=12;
					out<=141;
				end
				if(in == 550) begin
					state<=12;
					out<=142;
				end
				if(in == 551) begin
					state<=9;
					out<=143;
				end
				if(in == 552) begin
					state<=9;
					out<=144;
				end
				if(in == 553) begin
					state<=12;
					out<=145;
				end
				if(in == 554) begin
					state<=12;
					out<=146;
				end
				if(in == 555) begin
					state<=9;
					out<=147;
				end
				if(in == 556) begin
					state<=9;
					out<=148;
				end
				if(in == 557) begin
					state<=12;
					out<=149;
				end
				if(in == 558) begin
					state<=12;
					out<=150;
				end
				if(in == 559) begin
					state<=9;
					out<=151;
				end
				if(in == 560) begin
					state<=9;
					out<=152;
				end
				if(in == 561) begin
					state<=12;
					out<=153;
				end
				if(in == 562) begin
					state<=12;
					out<=154;
				end
				if(in == 563) begin
					state<=9;
					out<=155;
				end
				if(in == 564) begin
					state<=9;
					out<=156;
				end
				if(in == 565) begin
					state<=12;
					out<=157;
				end
				if(in == 566) begin
					state<=12;
					out<=158;
				end
				if(in == 567) begin
					state<=9;
					out<=159;
				end
				if(in == 568) begin
					state<=9;
					out<=160;
				end
				if(in == 569) begin
					state<=2;
					out<=161;
				end
				if(in == 570) begin
					state<=2;
					out<=162;
				end
				if(in == 571) begin
					state<=2;
					out<=163;
				end
				if(in == 572) begin
					state<=2;
					out<=164;
				end
				if(in == 573) begin
					state<=2;
					out<=165;
				end
				if(in == 574) begin
					state<=2;
					out<=166;
				end
				if(in == 575) begin
					state<=2;
					out<=167;
				end
				if(in == 576) begin
					state<=2;
					out<=168;
				end
				if(in == 577) begin
					state<=2;
					out<=169;
				end
				if(in == 578) begin
					state<=2;
					out<=170;
				end
				if(in == 579) begin
					state<=2;
					out<=171;
				end
				if(in == 580) begin
					state<=2;
					out<=172;
				end
				if(in == 581) begin
					state<=3;
					out<=173;
				end
				if(in == 582) begin
					state<=8;
					out<=174;
				end
				if(in == 583) begin
					state<=3;
					out<=175;
				end
				if(in == 584) begin
					state<=12;
					out<=176;
				end
				if(in == 585) begin
					state<=3;
					out<=177;
				end
				if(in == 586) begin
					state<=12;
					out<=178;
				end
				if(in == 587) begin
					state<=9;
					out<=179;
				end
				if(in == 588) begin
					state<=9;
					out<=180;
				end
				if(in == 589) begin
					state<=12;
					out<=181;
				end
				if(in == 590) begin
					state<=12;
					out<=182;
				end
				if(in == 591) begin
					state<=9;
					out<=183;
				end
				if(in == 592) begin
					state<=9;
					out<=184;
				end
				if(in == 593) begin
					state<=12;
					out<=185;
				end
				if(in == 594) begin
					state<=12;
					out<=186;
				end
				if(in == 595) begin
					state<=9;
					out<=187;
				end
				if(in == 596) begin
					state<=9;
					out<=188;
				end
				if(in == 597) begin
					state<=12;
					out<=189;
				end
				if(in == 598) begin
					state<=12;
					out<=190;
				end
				if(in == 599) begin
					state<=9;
					out<=191;
				end
				if(in == 600) begin
					state<=9;
					out<=192;
				end
				if(in == 601) begin
					state<=12;
					out<=193;
				end
				if(in == 602) begin
					state<=12;
					out<=194;
				end
				if(in == 603) begin
					state<=9;
					out<=195;
				end
				if(in == 604) begin
					state<=9;
					out<=196;
				end
				if(in == 605) begin
					state<=12;
					out<=197;
				end
				if(in == 606) begin
					state<=12;
					out<=198;
				end
				if(in == 607) begin
					state<=9;
					out<=199;
				end
				if(in == 608) begin
					state<=9;
					out<=200;
				end
				if(in == 609) begin
					state<=12;
					out<=201;
				end
				if(in == 610) begin
					state<=12;
					out<=202;
				end
				if(in == 611) begin
					state<=9;
					out<=203;
				end
				if(in == 612) begin
					state<=9;
					out<=204;
				end
				if(in == 613) begin
					state<=12;
					out<=205;
				end
				if(in == 614) begin
					state<=12;
					out<=206;
				end
				if(in == 615) begin
					state<=9;
					out<=207;
				end
				if(in == 616) begin
					state<=9;
					out<=208;
				end
				if(in == 617) begin
					state<=12;
					out<=209;
				end
				if(in == 618) begin
					state<=12;
					out<=210;
				end
				if(in == 619) begin
					state<=9;
					out<=211;
				end
				if(in == 620) begin
					state<=9;
					out<=212;
				end
				if(in == 621) begin
					state<=12;
					out<=213;
				end
				if(in == 622) begin
					state<=12;
					out<=214;
				end
				if(in == 623) begin
					state<=9;
					out<=215;
				end
				if(in == 624) begin
					state<=9;
					out<=216;
				end
				if(in == 625) begin
					state<=12;
					out<=217;
				end
				if(in == 626) begin
					state<=12;
					out<=218;
				end
				if(in == 627) begin
					state<=9;
					out<=219;
				end
				if(in == 628) begin
					state<=9;
					out<=220;
				end
				if(in == 629) begin
					state<=12;
					out<=221;
				end
				if(in == 630) begin
					state<=12;
					out<=222;
				end
				if(in == 631) begin
					state<=9;
					out<=223;
				end
				if(in == 632) begin
					state<=9;
					out<=224;
				end
				if(in == 633) begin
					state<=3;
					out<=225;
				end
				if(in == 634) begin
					state<=8;
					out<=226;
				end
				if(in == 635) begin
					state<=3;
					out<=227;
				end
				if(in == 636) begin
					state<=12;
					out<=228;
				end
				if(in == 637) begin
					state<=3;
					out<=229;
				end
				if(in == 638) begin
					state<=12;
					out<=230;
				end
				if(in == 639) begin
					state<=9;
					out<=231;
				end
				if(in == 640) begin
					state<=9;
					out<=232;
				end
				if(in == 641) begin
					state<=12;
					out<=233;
				end
				if(in == 642) begin
					state<=12;
					out<=234;
				end
				if(in == 643) begin
					state<=9;
					out<=235;
				end
				if(in == 644) begin
					state<=9;
					out<=236;
				end
				if(in == 645) begin
					state<=12;
					out<=237;
				end
				if(in == 646) begin
					state<=12;
					out<=238;
				end
				if(in == 647) begin
					state<=9;
					out<=239;
				end
				if(in == 648) begin
					state<=9;
					out<=240;
				end
				if(in == 649) begin
					state<=12;
					out<=241;
				end
				if(in == 650) begin
					state<=12;
					out<=242;
				end
				if(in == 651) begin
					state<=9;
					out<=243;
				end
				if(in == 652) begin
					state<=9;
					out<=244;
				end
				if(in == 653) begin
					state<=12;
					out<=245;
				end
				if(in == 654) begin
					state<=12;
					out<=246;
				end
				if(in == 655) begin
					state<=9;
					out<=247;
				end
				if(in == 656) begin
					state<=9;
					out<=248;
				end
				if(in == 657) begin
					state<=12;
					out<=249;
				end
				if(in == 658) begin
					state<=12;
					out<=250;
				end
				if(in == 659) begin
					state<=9;
					out<=251;
				end
				if(in == 660) begin
					state<=9;
					out<=252;
				end
				if(in == 661) begin
					state<=12;
					out<=253;
				end
				if(in == 662) begin
					state<=12;
					out<=254;
				end
				if(in == 663) begin
					state<=9;
					out<=255;
				end
				if(in == 664) begin
					state<=9;
					out<=0;
				end
				if(in == 665) begin
					state<=12;
					out<=1;
				end
				if(in == 666) begin
					state<=12;
					out<=2;
				end
				if(in == 667) begin
					state<=9;
					out<=3;
				end
				if(in == 668) begin
					state<=9;
					out<=4;
				end
				if(in == 669) begin
					state<=12;
					out<=5;
				end
				if(in == 670) begin
					state<=12;
					out<=6;
				end
				if(in == 671) begin
					state<=9;
					out<=7;
				end
				if(in == 672) begin
					state<=9;
					out<=8;
				end
				if(in == 673) begin
					state<=12;
					out<=9;
				end
				if(in == 674) begin
					state<=12;
					out<=10;
				end
				if(in == 675) begin
					state<=9;
					out<=11;
				end
				if(in == 676) begin
					state<=9;
					out<=12;
				end
				if(in == 677) begin
					state<=12;
					out<=13;
				end
				if(in == 678) begin
					state<=12;
					out<=14;
				end
				if(in == 679) begin
					state<=9;
					out<=15;
				end
				if(in == 680) begin
					state<=9;
					out<=16;
				end
				if(in == 681) begin
					state<=12;
					out<=17;
				end
				if(in == 682) begin
					state<=12;
					out<=18;
				end
				if(in == 683) begin
					state<=9;
					out<=19;
				end
				if(in == 684) begin
					state<=9;
					out<=20;
				end
				if(in == 685) begin
					state<=2;
					out<=21;
				end
				if(in == 686) begin
					state<=2;
					out<=22;
				end
				if(in == 687) begin
					state<=2;
					out<=23;
				end
				if(in == 688) begin
					state<=2;
					out<=24;
				end
				if(in == 689) begin
					state<=2;
					out<=25;
				end
				if(in == 690) begin
					state<=2;
					out<=26;
				end
				if(in == 691) begin
					state<=2;
					out<=27;
				end
				if(in == 692) begin
					state<=2;
					out<=28;
				end
				if(in == 693) begin
					state<=2;
					out<=29;
				end
				if(in == 694) begin
					state<=2;
					out<=30;
				end
				if(in == 695) begin
					state<=2;
					out<=31;
				end
				if(in == 696) begin
					state<=2;
					out<=32;
				end
				if(in == 697) begin
					state<=3;
					out<=33;
				end
				if(in == 698) begin
					state<=8;
					out<=34;
				end
				if(in == 699) begin
					state<=3;
					out<=35;
				end
				if(in == 700) begin
					state<=12;
					out<=36;
				end
				if(in == 701) begin
					state<=3;
					out<=37;
				end
				if(in == 702) begin
					state<=12;
					out<=38;
				end
				if(in == 703) begin
					state<=9;
					out<=39;
				end
				if(in == 704) begin
					state<=9;
					out<=40;
				end
				if(in == 705) begin
					state<=12;
					out<=41;
				end
				if(in == 706) begin
					state<=12;
					out<=42;
				end
				if(in == 707) begin
					state<=9;
					out<=43;
				end
				if(in == 708) begin
					state<=9;
					out<=44;
				end
				if(in == 709) begin
					state<=12;
					out<=45;
				end
				if(in == 710) begin
					state<=12;
					out<=46;
				end
				if(in == 711) begin
					state<=9;
					out<=47;
				end
				if(in == 712) begin
					state<=9;
					out<=48;
				end
				if(in == 713) begin
					state<=12;
					out<=49;
				end
				if(in == 714) begin
					state<=12;
					out<=50;
				end
				if(in == 715) begin
					state<=9;
					out<=51;
				end
				if(in == 716) begin
					state<=9;
					out<=52;
				end
				if(in == 717) begin
					state<=12;
					out<=53;
				end
				if(in == 718) begin
					state<=12;
					out<=54;
				end
				if(in == 719) begin
					state<=9;
					out<=55;
				end
				if(in == 720) begin
					state<=9;
					out<=56;
				end
				if(in == 721) begin
					state<=12;
					out<=57;
				end
				if(in == 722) begin
					state<=12;
					out<=58;
				end
				if(in == 723) begin
					state<=9;
					out<=59;
				end
				if(in == 724) begin
					state<=9;
					out<=60;
				end
				if(in == 725) begin
					state<=12;
					out<=61;
				end
				if(in == 726) begin
					state<=12;
					out<=62;
				end
				if(in == 727) begin
					state<=9;
					out<=63;
				end
				if(in == 728) begin
					state<=9;
					out<=64;
				end
				if(in == 729) begin
					state<=12;
					out<=65;
				end
				if(in == 730) begin
					state<=12;
					out<=66;
				end
				if(in == 731) begin
					state<=9;
					out<=67;
				end
				if(in == 732) begin
					state<=9;
					out<=68;
				end
				if(in == 733) begin
					state<=12;
					out<=69;
				end
				if(in == 734) begin
					state<=12;
					out<=70;
				end
				if(in == 735) begin
					state<=9;
					out<=71;
				end
				if(in == 736) begin
					state<=9;
					out<=72;
				end
				if(in == 737) begin
					state<=12;
					out<=73;
				end
				if(in == 738) begin
					state<=12;
					out<=74;
				end
				if(in == 739) begin
					state<=9;
					out<=75;
				end
				if(in == 740) begin
					state<=9;
					out<=76;
				end
				if(in == 741) begin
					state<=12;
					out<=77;
				end
				if(in == 742) begin
					state<=12;
					out<=78;
				end
				if(in == 743) begin
					state<=9;
					out<=79;
				end
				if(in == 744) begin
					state<=9;
					out<=80;
				end
				if(in == 745) begin
					state<=12;
					out<=81;
				end
				if(in == 746) begin
					state<=12;
					out<=82;
				end
				if(in == 747) begin
					state<=9;
					out<=83;
				end
				if(in == 748) begin
					state<=9;
					out<=84;
				end
				if(in == 749) begin
					state<=3;
					out<=85;
				end
				if(in == 750) begin
					state<=8;
					out<=86;
				end
				if(in == 751) begin
					state<=3;
					out<=87;
				end
				if(in == 752) begin
					state<=12;
					out<=88;
				end
				if(in == 753) begin
					state<=3;
					out<=89;
				end
				if(in == 754) begin
					state<=12;
					out<=90;
				end
				if(in == 755) begin
					state<=9;
					out<=91;
				end
				if(in == 756) begin
					state<=9;
					out<=92;
				end
				if(in == 757) begin
					state<=12;
					out<=93;
				end
				if(in == 758) begin
					state<=12;
					out<=94;
				end
				if(in == 759) begin
					state<=9;
					out<=95;
				end
				if(in == 760) begin
					state<=9;
					out<=96;
				end
				if(in == 761) begin
					state<=12;
					out<=97;
				end
				if(in == 762) begin
					state<=12;
					out<=98;
				end
				if(in == 763) begin
					state<=9;
					out<=99;
				end
				if(in == 764) begin
					state<=9;
					out<=100;
				end
				if(in == 765) begin
					state<=12;
					out<=101;
				end
				if(in == 766) begin
					state<=12;
					out<=102;
				end
				if(in == 767) begin
					state<=9;
					out<=103;
				end
				if(in == 768) begin
					state<=9;
					out<=104;
				end
				if(in == 769) begin
					state<=12;
					out<=105;
				end
				if(in == 770) begin
					state<=12;
					out<=106;
				end
				if(in == 771) begin
					state<=9;
					out<=107;
				end
				if(in == 772) begin
					state<=9;
					out<=108;
				end
				if(in == 773) begin
					state<=12;
					out<=109;
				end
				if(in == 774) begin
					state<=12;
					out<=110;
				end
				if(in == 775) begin
					state<=9;
					out<=111;
				end
				if(in == 776) begin
					state<=9;
					out<=112;
				end
				if(in == 777) begin
					state<=12;
					out<=113;
				end
				if(in == 778) begin
					state<=12;
					out<=114;
				end
				if(in == 779) begin
					state<=9;
					out<=115;
				end
				if(in == 780) begin
					state<=9;
					out<=116;
				end
				if(in == 781) begin
					state<=12;
					out<=117;
				end
				if(in == 782) begin
					state<=12;
					out<=118;
				end
				if(in == 783) begin
					state<=9;
					out<=119;
				end
				if(in == 784) begin
					state<=9;
					out<=120;
				end
				if(in == 785) begin
					state<=12;
					out<=121;
				end
				if(in == 786) begin
					state<=12;
					out<=122;
				end
				if(in == 787) begin
					state<=9;
					out<=123;
				end
				if(in == 788) begin
					state<=9;
					out<=124;
				end
				if(in == 789) begin
					state<=12;
					out<=125;
				end
				if(in == 790) begin
					state<=12;
					out<=126;
				end
				if(in == 791) begin
					state<=9;
					out<=127;
				end
				if(in == 792) begin
					state<=9;
					out<=128;
				end
				if(in == 793) begin
					state<=12;
					out<=129;
				end
				if(in == 794) begin
					state<=12;
					out<=130;
				end
				if(in == 795) begin
					state<=9;
					out<=131;
				end
				if(in == 796) begin
					state<=9;
					out<=132;
				end
				if(in == 797) begin
					state<=12;
					out<=133;
				end
				if(in == 798) begin
					state<=12;
					out<=134;
				end
				if(in == 799) begin
					state<=9;
					out<=135;
				end
				if(in == 800) begin
					state<=9;
					out<=136;
				end
				if(in == 801) begin
					state<=2;
					out<=137;
				end
				if(in == 802) begin
					state<=2;
					out<=138;
				end
				if(in == 803) begin
					state<=2;
					out<=139;
				end
				if(in == 804) begin
					state<=2;
					out<=140;
				end
				if(in == 805) begin
					state<=2;
					out<=141;
				end
				if(in == 806) begin
					state<=2;
					out<=142;
				end
				if(in == 807) begin
					state<=2;
					out<=143;
				end
				if(in == 808) begin
					state<=2;
					out<=144;
				end
				if(in == 809) begin
					state<=2;
					out<=145;
				end
				if(in == 810) begin
					state<=2;
					out<=146;
				end
				if(in == 811) begin
					state<=2;
					out<=147;
				end
				if(in == 812) begin
					state<=2;
					out<=148;
				end
				if(in == 813) begin
					state<=3;
					out<=149;
				end
				if(in == 814) begin
					state<=8;
					out<=150;
				end
				if(in == 815) begin
					state<=3;
					out<=151;
				end
				if(in == 816) begin
					state<=12;
					out<=152;
				end
				if(in == 817) begin
					state<=3;
					out<=153;
				end
				if(in == 818) begin
					state<=12;
					out<=154;
				end
				if(in == 819) begin
					state<=9;
					out<=155;
				end
				if(in == 820) begin
					state<=9;
					out<=156;
				end
				if(in == 821) begin
					state<=12;
					out<=157;
				end
				if(in == 822) begin
					state<=12;
					out<=158;
				end
				if(in == 823) begin
					state<=9;
					out<=159;
				end
				if(in == 824) begin
					state<=9;
					out<=160;
				end
				if(in == 825) begin
					state<=12;
					out<=161;
				end
				if(in == 826) begin
					state<=12;
					out<=162;
				end
				if(in == 827) begin
					state<=9;
					out<=163;
				end
				if(in == 828) begin
					state<=9;
					out<=164;
				end
				if(in == 829) begin
					state<=12;
					out<=165;
				end
				if(in == 830) begin
					state<=12;
					out<=166;
				end
				if(in == 831) begin
					state<=9;
					out<=167;
				end
				if(in == 832) begin
					state<=9;
					out<=168;
				end
				if(in == 833) begin
					state<=12;
					out<=169;
				end
				if(in == 834) begin
					state<=12;
					out<=170;
				end
				if(in == 835) begin
					state<=9;
					out<=171;
				end
				if(in == 836) begin
					state<=9;
					out<=172;
				end
				if(in == 837) begin
					state<=12;
					out<=173;
				end
				if(in == 838) begin
					state<=12;
					out<=174;
				end
				if(in == 839) begin
					state<=9;
					out<=175;
				end
				if(in == 840) begin
					state<=9;
					out<=176;
				end
				if(in == 841) begin
					state<=12;
					out<=177;
				end
				if(in == 842) begin
					state<=12;
					out<=178;
				end
				if(in == 843) begin
					state<=9;
					out<=179;
				end
				if(in == 844) begin
					state<=9;
					out<=180;
				end
				if(in == 845) begin
					state<=12;
					out<=181;
				end
				if(in == 846) begin
					state<=12;
					out<=182;
				end
				if(in == 847) begin
					state<=9;
					out<=183;
				end
				if(in == 848) begin
					state<=9;
					out<=184;
				end
				if(in == 849) begin
					state<=12;
					out<=185;
				end
				if(in == 850) begin
					state<=12;
					out<=186;
				end
				if(in == 851) begin
					state<=9;
					out<=187;
				end
				if(in == 852) begin
					state<=9;
					out<=188;
				end
				if(in == 853) begin
					state<=12;
					out<=189;
				end
				if(in == 854) begin
					state<=12;
					out<=190;
				end
				if(in == 855) begin
					state<=9;
					out<=191;
				end
				if(in == 856) begin
					state<=9;
					out<=192;
				end
				if(in == 857) begin
					state<=12;
					out<=193;
				end
				if(in == 858) begin
					state<=12;
					out<=194;
				end
				if(in == 859) begin
					state<=9;
					out<=195;
				end
				if(in == 860) begin
					state<=9;
					out<=196;
				end
				if(in == 861) begin
					state<=12;
					out<=197;
				end
				if(in == 862) begin
					state<=12;
					out<=198;
				end
				if(in == 863) begin
					state<=9;
					out<=199;
				end
				if(in == 864) begin
					state<=9;
					out<=200;
				end
				if(in == 865) begin
					state<=3;
					out<=201;
				end
				if(in == 866) begin
					state<=8;
					out<=202;
				end
				if(in == 867) begin
					state<=3;
					out<=203;
				end
				if(in == 868) begin
					state<=12;
					out<=204;
				end
				if(in == 869) begin
					state<=3;
					out<=205;
				end
				if(in == 870) begin
					state<=12;
					out<=206;
				end
				if(in == 871) begin
					state<=9;
					out<=207;
				end
				if(in == 872) begin
					state<=9;
					out<=208;
				end
				if(in == 873) begin
					state<=12;
					out<=209;
				end
				if(in == 874) begin
					state<=12;
					out<=210;
				end
				if(in == 875) begin
					state<=9;
					out<=211;
				end
				if(in == 876) begin
					state<=9;
					out<=212;
				end
				if(in == 877) begin
					state<=12;
					out<=213;
				end
				if(in == 878) begin
					state<=12;
					out<=214;
				end
				if(in == 879) begin
					state<=9;
					out<=215;
				end
				if(in == 880) begin
					state<=9;
					out<=216;
				end
				if(in == 881) begin
					state<=12;
					out<=217;
				end
				if(in == 882) begin
					state<=12;
					out<=218;
				end
				if(in == 883) begin
					state<=9;
					out<=219;
				end
				if(in == 884) begin
					state<=9;
					out<=220;
				end
				if(in == 885) begin
					state<=12;
					out<=221;
				end
				if(in == 886) begin
					state<=12;
					out<=222;
				end
				if(in == 887) begin
					state<=9;
					out<=223;
				end
				if(in == 888) begin
					state<=9;
					out<=224;
				end
				if(in == 889) begin
					state<=12;
					out<=225;
				end
				if(in == 890) begin
					state<=12;
					out<=226;
				end
				if(in == 891) begin
					state<=9;
					out<=227;
				end
				if(in == 892) begin
					state<=9;
					out<=228;
				end
				if(in == 893) begin
					state<=12;
					out<=229;
				end
				if(in == 894) begin
					state<=12;
					out<=230;
				end
				if(in == 895) begin
					state<=9;
					out<=231;
				end
				if(in == 896) begin
					state<=9;
					out<=232;
				end
				if(in == 897) begin
					state<=12;
					out<=233;
				end
				if(in == 898) begin
					state<=12;
					out<=234;
				end
				if(in == 899) begin
					state<=9;
					out<=235;
				end
				if(in == 900) begin
					state<=9;
					out<=236;
				end
				if(in == 901) begin
					state<=12;
					out<=237;
				end
				if(in == 902) begin
					state<=12;
					out<=238;
				end
				if(in == 903) begin
					state<=9;
					out<=239;
				end
				if(in == 904) begin
					state<=9;
					out<=240;
				end
				if(in == 905) begin
					state<=12;
					out<=241;
				end
				if(in == 906) begin
					state<=12;
					out<=242;
				end
				if(in == 907) begin
					state<=9;
					out<=243;
				end
				if(in == 908) begin
					state<=9;
					out<=244;
				end
				if(in == 909) begin
					state<=12;
					out<=245;
				end
				if(in == 910) begin
					state<=12;
					out<=246;
				end
				if(in == 911) begin
					state<=9;
					out<=247;
				end
				if(in == 912) begin
					state<=9;
					out<=248;
				end
				if(in == 913) begin
					state<=12;
					out<=249;
				end
				if(in == 914) begin
					state<=12;
					out<=250;
				end
				if(in == 915) begin
					state<=9;
					out<=251;
				end
				if(in == 916) begin
					state<=9;
					out<=252;
				end
				if(in == 917) begin
					state<=2;
					out<=253;
				end
				if(in == 918) begin
					state<=2;
					out<=254;
				end
				if(in == 919) begin
					state<=2;
					out<=255;
				end
				if(in == 920) begin
					state<=2;
					out<=0;
				end
				if(in == 921) begin
					state<=2;
					out<=1;
				end
				if(in == 922) begin
					state<=2;
					out<=2;
				end
				if(in == 923) begin
					state<=2;
					out<=3;
				end
				if(in == 924) begin
					state<=2;
					out<=4;
				end
				if(in == 925) begin
					state<=2;
					out<=5;
				end
				if(in == 926) begin
					state<=2;
					out<=6;
				end
				if(in == 927) begin
					state<=2;
					out<=7;
				end
				if(in == 928) begin
					state<=2;
					out<=8;
				end
			end
			9: begin
				if(in == 0) begin
					state<=3;
					out<=9;
				end
				if(in == 1) begin
					state<=1;
					out<=10;
				end
				if(in == 2) begin
					state<=9;
					out<=11;
				end
				if(in == 3) begin
					state<=3;
					out<=12;
				end
				if(in == 4) begin
					state<=10;
					out<=13;
				end
				if(in == 5) begin
					state<=3;
					out<=14;
				end
				if(in == 6) begin
					state<=10;
					out<=15;
				end
				if(in == 7) begin
					state<=10;
					out<=16;
				end
				if(in == 8) begin
					state<=10;
					out<=17;
				end
				if(in == 9) begin
					state<=10;
					out<=18;
				end
				if(in == 10) begin
					state<=10;
					out<=19;
				end
				if(in == 11) begin
					state<=10;
					out<=20;
				end
				if(in == 12) begin
					state<=10;
					out<=21;
				end
				if(in == 13) begin
					state<=10;
					out<=22;
				end
				if(in == 14) begin
					state<=10;
					out<=23;
				end
				if(in == 15) begin
					state<=10;
					out<=24;
				end
				if(in == 16) begin
					state<=10;
					out<=25;
				end
				if(in == 17) begin
					state<=10;
					out<=26;
				end
				if(in == 18) begin
					state<=10;
					out<=27;
				end
				if(in == 19) begin
					state<=10;
					out<=28;
				end
				if(in == 20) begin
					state<=10;
					out<=29;
				end
				if(in == 21) begin
					state<=10;
					out<=30;
				end
				if(in == 22) begin
					state<=10;
					out<=31;
				end
				if(in == 23) begin
					state<=10;
					out<=32;
				end
				if(in == 24) begin
					state<=10;
					out<=33;
				end
				if(in == 25) begin
					state<=10;
					out<=34;
				end
				if(in == 26) begin
					state<=10;
					out<=35;
				end
				if(in == 27) begin
					state<=10;
					out<=36;
				end
				if(in == 28) begin
					state<=10;
					out<=37;
				end
				if(in == 29) begin
					state<=10;
					out<=38;
				end
				if(in == 30) begin
					state<=10;
					out<=39;
				end
				if(in == 31) begin
					state<=10;
					out<=40;
				end
				if(in == 32) begin
					state<=10;
					out<=41;
				end
				if(in == 33) begin
					state<=10;
					out<=42;
				end
				if(in == 34) begin
					state<=10;
					out<=43;
				end
				if(in == 35) begin
					state<=10;
					out<=44;
				end
				if(in == 36) begin
					state<=10;
					out<=45;
				end
				if(in == 37) begin
					state<=10;
					out<=46;
				end
				if(in == 38) begin
					state<=10;
					out<=47;
				end
				if(in == 39) begin
					state<=10;
					out<=48;
				end
				if(in == 40) begin
					state<=10;
					out<=49;
				end
				if(in == 41) begin
					state<=10;
					out<=50;
				end
				if(in == 42) begin
					state<=10;
					out<=51;
				end
				if(in == 43) begin
					state<=10;
					out<=52;
				end
				if(in == 44) begin
					state<=10;
					out<=53;
				end
				if(in == 45) begin
					state<=10;
					out<=54;
				end
				if(in == 46) begin
					state<=10;
					out<=55;
				end
				if(in == 47) begin
					state<=10;
					out<=56;
				end
				if(in == 48) begin
					state<=10;
					out<=57;
				end
				if(in == 49) begin
					state<=10;
					out<=58;
				end
				if(in == 50) begin
					state<=10;
					out<=59;
				end
				if(in == 51) begin
					state<=10;
					out<=60;
				end
				if(in == 52) begin
					state<=10;
					out<=61;
				end
				if(in == 53) begin
					state<=3;
					out<=62;
				end
				if(in == 54) begin
					state<=9;
					out<=63;
				end
				if(in == 55) begin
					state<=3;
					out<=64;
				end
				if(in == 56) begin
					state<=10;
					out<=65;
				end
				if(in == 57) begin
					state<=3;
					out<=66;
				end
				if(in == 58) begin
					state<=10;
					out<=67;
				end
				if(in == 59) begin
					state<=10;
					out<=68;
				end
				if(in == 60) begin
					state<=10;
					out<=69;
				end
				if(in == 61) begin
					state<=10;
					out<=70;
				end
				if(in == 62) begin
					state<=10;
					out<=71;
				end
				if(in == 63) begin
					state<=10;
					out<=72;
				end
				if(in == 64) begin
					state<=10;
					out<=73;
				end
				if(in == 65) begin
					state<=10;
					out<=74;
				end
				if(in == 66) begin
					state<=10;
					out<=75;
				end
				if(in == 67) begin
					state<=10;
					out<=76;
				end
				if(in == 68) begin
					state<=10;
					out<=77;
				end
				if(in == 69) begin
					state<=10;
					out<=78;
				end
				if(in == 70) begin
					state<=10;
					out<=79;
				end
				if(in == 71) begin
					state<=10;
					out<=80;
				end
				if(in == 72) begin
					state<=10;
					out<=81;
				end
				if(in == 73) begin
					state<=10;
					out<=82;
				end
				if(in == 74) begin
					state<=10;
					out<=83;
				end
				if(in == 75) begin
					state<=10;
					out<=84;
				end
				if(in == 76) begin
					state<=10;
					out<=85;
				end
				if(in == 77) begin
					state<=10;
					out<=86;
				end
				if(in == 78) begin
					state<=10;
					out<=87;
				end
				if(in == 79) begin
					state<=10;
					out<=88;
				end
				if(in == 80) begin
					state<=10;
					out<=89;
				end
				if(in == 81) begin
					state<=10;
					out<=90;
				end
				if(in == 82) begin
					state<=10;
					out<=91;
				end
				if(in == 83) begin
					state<=10;
					out<=92;
				end
				if(in == 84) begin
					state<=10;
					out<=93;
				end
				if(in == 85) begin
					state<=10;
					out<=94;
				end
				if(in == 86) begin
					state<=10;
					out<=95;
				end
				if(in == 87) begin
					state<=10;
					out<=96;
				end
				if(in == 88) begin
					state<=10;
					out<=97;
				end
				if(in == 89) begin
					state<=10;
					out<=98;
				end
				if(in == 90) begin
					state<=10;
					out<=99;
				end
				if(in == 91) begin
					state<=10;
					out<=100;
				end
				if(in == 92) begin
					state<=10;
					out<=101;
				end
				if(in == 93) begin
					state<=10;
					out<=102;
				end
				if(in == 94) begin
					state<=10;
					out<=103;
				end
				if(in == 95) begin
					state<=10;
					out<=104;
				end
				if(in == 96) begin
					state<=10;
					out<=105;
				end
				if(in == 97) begin
					state<=10;
					out<=106;
				end
				if(in == 98) begin
					state<=10;
					out<=107;
				end
				if(in == 99) begin
					state<=10;
					out<=108;
				end
				if(in == 100) begin
					state<=10;
					out<=109;
				end
				if(in == 101) begin
					state<=10;
					out<=110;
				end
				if(in == 102) begin
					state<=10;
					out<=111;
				end
				if(in == 103) begin
					state<=10;
					out<=112;
				end
				if(in == 104) begin
					state<=10;
					out<=113;
				end
				if(in == 105) begin
					state<=2;
					out<=114;
				end
				if(in == 106) begin
					state<=2;
					out<=115;
				end
				if(in == 107) begin
					state<=2;
					out<=116;
				end
				if(in == 108) begin
					state<=2;
					out<=117;
				end
				if(in == 109) begin
					state<=2;
					out<=118;
				end
				if(in == 110) begin
					state<=2;
					out<=119;
				end
				if(in == 111) begin
					state<=2;
					out<=120;
				end
				if(in == 112) begin
					state<=2;
					out<=121;
				end
				if(in == 113) begin
					state<=2;
					out<=122;
				end
				if(in == 114) begin
					state<=2;
					out<=123;
				end
				if(in == 115) begin
					state<=2;
					out<=124;
				end
				if(in == 116) begin
					state<=2;
					out<=125;
				end
				if(in == 117) begin
					state<=3;
					out<=126;
				end
				if(in == 118) begin
					state<=9;
					out<=127;
				end
				if(in == 119) begin
					state<=3;
					out<=128;
				end
				if(in == 120) begin
					state<=10;
					out<=129;
				end
				if(in == 121) begin
					state<=3;
					out<=130;
				end
				if(in == 122) begin
					state<=10;
					out<=131;
				end
				if(in == 123) begin
					state<=10;
					out<=132;
				end
				if(in == 124) begin
					state<=10;
					out<=133;
				end
				if(in == 125) begin
					state<=10;
					out<=134;
				end
				if(in == 126) begin
					state<=10;
					out<=135;
				end
				if(in == 127) begin
					state<=10;
					out<=136;
				end
				if(in == 128) begin
					state<=10;
					out<=137;
				end
				if(in == 129) begin
					state<=10;
					out<=138;
				end
				if(in == 130) begin
					state<=10;
					out<=139;
				end
				if(in == 131) begin
					state<=10;
					out<=140;
				end
				if(in == 132) begin
					state<=10;
					out<=141;
				end
				if(in == 133) begin
					state<=10;
					out<=142;
				end
				if(in == 134) begin
					state<=10;
					out<=143;
				end
				if(in == 135) begin
					state<=10;
					out<=144;
				end
				if(in == 136) begin
					state<=10;
					out<=145;
				end
				if(in == 137) begin
					state<=10;
					out<=146;
				end
				if(in == 138) begin
					state<=10;
					out<=147;
				end
				if(in == 139) begin
					state<=10;
					out<=148;
				end
				if(in == 140) begin
					state<=10;
					out<=149;
				end
				if(in == 141) begin
					state<=10;
					out<=150;
				end
				if(in == 142) begin
					state<=10;
					out<=151;
				end
				if(in == 143) begin
					state<=10;
					out<=152;
				end
				if(in == 144) begin
					state<=10;
					out<=153;
				end
				if(in == 145) begin
					state<=10;
					out<=154;
				end
				if(in == 146) begin
					state<=10;
					out<=155;
				end
				if(in == 147) begin
					state<=10;
					out<=156;
				end
				if(in == 148) begin
					state<=10;
					out<=157;
				end
				if(in == 149) begin
					state<=10;
					out<=158;
				end
				if(in == 150) begin
					state<=10;
					out<=159;
				end
				if(in == 151) begin
					state<=10;
					out<=160;
				end
				if(in == 152) begin
					state<=10;
					out<=161;
				end
				if(in == 153) begin
					state<=10;
					out<=162;
				end
				if(in == 154) begin
					state<=10;
					out<=163;
				end
				if(in == 155) begin
					state<=10;
					out<=164;
				end
				if(in == 156) begin
					state<=10;
					out<=165;
				end
				if(in == 157) begin
					state<=10;
					out<=166;
				end
				if(in == 158) begin
					state<=10;
					out<=167;
				end
				if(in == 159) begin
					state<=10;
					out<=168;
				end
				if(in == 160) begin
					state<=10;
					out<=169;
				end
				if(in == 161) begin
					state<=10;
					out<=170;
				end
				if(in == 162) begin
					state<=10;
					out<=171;
				end
				if(in == 163) begin
					state<=10;
					out<=172;
				end
				if(in == 164) begin
					state<=10;
					out<=173;
				end
				if(in == 165) begin
					state<=10;
					out<=174;
				end
				if(in == 166) begin
					state<=10;
					out<=175;
				end
				if(in == 167) begin
					state<=10;
					out<=176;
				end
				if(in == 168) begin
					state<=10;
					out<=177;
				end
				if(in == 169) begin
					state<=3;
					out<=178;
				end
				if(in == 170) begin
					state<=9;
					out<=179;
				end
				if(in == 171) begin
					state<=3;
					out<=180;
				end
				if(in == 172) begin
					state<=10;
					out<=181;
				end
				if(in == 173) begin
					state<=3;
					out<=182;
				end
				if(in == 174) begin
					state<=10;
					out<=183;
				end
				if(in == 175) begin
					state<=10;
					out<=184;
				end
				if(in == 176) begin
					state<=10;
					out<=185;
				end
				if(in == 177) begin
					state<=10;
					out<=186;
				end
				if(in == 178) begin
					state<=10;
					out<=187;
				end
				if(in == 179) begin
					state<=10;
					out<=188;
				end
				if(in == 180) begin
					state<=10;
					out<=189;
				end
				if(in == 181) begin
					state<=10;
					out<=190;
				end
				if(in == 182) begin
					state<=10;
					out<=191;
				end
				if(in == 183) begin
					state<=10;
					out<=192;
				end
				if(in == 184) begin
					state<=10;
					out<=193;
				end
				if(in == 185) begin
					state<=10;
					out<=194;
				end
				if(in == 186) begin
					state<=10;
					out<=195;
				end
				if(in == 187) begin
					state<=10;
					out<=196;
				end
				if(in == 188) begin
					state<=10;
					out<=197;
				end
				if(in == 189) begin
					state<=10;
					out<=198;
				end
				if(in == 190) begin
					state<=10;
					out<=199;
				end
				if(in == 191) begin
					state<=10;
					out<=200;
				end
				if(in == 192) begin
					state<=10;
					out<=201;
				end
				if(in == 193) begin
					state<=10;
					out<=202;
				end
				if(in == 194) begin
					state<=10;
					out<=203;
				end
				if(in == 195) begin
					state<=10;
					out<=204;
				end
				if(in == 196) begin
					state<=10;
					out<=205;
				end
				if(in == 197) begin
					state<=10;
					out<=206;
				end
				if(in == 198) begin
					state<=10;
					out<=207;
				end
				if(in == 199) begin
					state<=10;
					out<=208;
				end
				if(in == 200) begin
					state<=10;
					out<=209;
				end
				if(in == 201) begin
					state<=10;
					out<=210;
				end
				if(in == 202) begin
					state<=10;
					out<=211;
				end
				if(in == 203) begin
					state<=10;
					out<=212;
				end
				if(in == 204) begin
					state<=10;
					out<=213;
				end
				if(in == 205) begin
					state<=10;
					out<=214;
				end
				if(in == 206) begin
					state<=10;
					out<=215;
				end
				if(in == 207) begin
					state<=10;
					out<=216;
				end
				if(in == 208) begin
					state<=10;
					out<=217;
				end
				if(in == 209) begin
					state<=10;
					out<=218;
				end
				if(in == 210) begin
					state<=10;
					out<=219;
				end
				if(in == 211) begin
					state<=10;
					out<=220;
				end
				if(in == 212) begin
					state<=10;
					out<=221;
				end
				if(in == 213) begin
					state<=10;
					out<=222;
				end
				if(in == 214) begin
					state<=10;
					out<=223;
				end
				if(in == 215) begin
					state<=10;
					out<=224;
				end
				if(in == 216) begin
					state<=10;
					out<=225;
				end
				if(in == 217) begin
					state<=10;
					out<=226;
				end
				if(in == 218) begin
					state<=10;
					out<=227;
				end
				if(in == 219) begin
					state<=10;
					out<=228;
				end
				if(in == 220) begin
					state<=10;
					out<=229;
				end
				if(in == 221) begin
					state<=2;
					out<=230;
				end
				if(in == 222) begin
					state<=2;
					out<=231;
				end
				if(in == 223) begin
					state<=2;
					out<=232;
				end
				if(in == 224) begin
					state<=2;
					out<=233;
				end
				if(in == 225) begin
					state<=2;
					out<=234;
				end
				if(in == 226) begin
					state<=2;
					out<=235;
				end
				if(in == 227) begin
					state<=2;
					out<=236;
				end
				if(in == 228) begin
					state<=2;
					out<=237;
				end
				if(in == 229) begin
					state<=2;
					out<=238;
				end
				if(in == 230) begin
					state<=2;
					out<=239;
				end
				if(in == 231) begin
					state<=2;
					out<=240;
				end
				if(in == 232) begin
					state<=2;
					out<=241;
				end
				if(in == 233) begin
					state<=3;
					out<=242;
				end
				if(in == 234) begin
					state<=9;
					out<=243;
				end
				if(in == 235) begin
					state<=3;
					out<=244;
				end
				if(in == 236) begin
					state<=10;
					out<=245;
				end
				if(in == 237) begin
					state<=3;
					out<=246;
				end
				if(in == 238) begin
					state<=10;
					out<=247;
				end
				if(in == 239) begin
					state<=10;
					out<=248;
				end
				if(in == 240) begin
					state<=10;
					out<=249;
				end
				if(in == 241) begin
					state<=10;
					out<=250;
				end
				if(in == 242) begin
					state<=10;
					out<=251;
				end
				if(in == 243) begin
					state<=10;
					out<=252;
				end
				if(in == 244) begin
					state<=10;
					out<=253;
				end
				if(in == 245) begin
					state<=10;
					out<=254;
				end
				if(in == 246) begin
					state<=10;
					out<=255;
				end
				if(in == 247) begin
					state<=10;
					out<=0;
				end
				if(in == 248) begin
					state<=10;
					out<=1;
				end
				if(in == 249) begin
					state<=10;
					out<=2;
				end
				if(in == 250) begin
					state<=10;
					out<=3;
				end
				if(in == 251) begin
					state<=10;
					out<=4;
				end
				if(in == 252) begin
					state<=10;
					out<=5;
				end
				if(in == 253) begin
					state<=10;
					out<=6;
				end
				if(in == 254) begin
					state<=10;
					out<=7;
				end
				if(in == 255) begin
					state<=10;
					out<=8;
				end
				if(in == 256) begin
					state<=10;
					out<=9;
				end
				if(in == 257) begin
					state<=10;
					out<=10;
				end
				if(in == 258) begin
					state<=10;
					out<=11;
				end
				if(in == 259) begin
					state<=10;
					out<=12;
				end
				if(in == 260) begin
					state<=10;
					out<=13;
				end
				if(in == 261) begin
					state<=10;
					out<=14;
				end
				if(in == 262) begin
					state<=10;
					out<=15;
				end
				if(in == 263) begin
					state<=10;
					out<=16;
				end
				if(in == 264) begin
					state<=10;
					out<=17;
				end
				if(in == 265) begin
					state<=10;
					out<=18;
				end
				if(in == 266) begin
					state<=10;
					out<=19;
				end
				if(in == 267) begin
					state<=10;
					out<=20;
				end
				if(in == 268) begin
					state<=10;
					out<=21;
				end
				if(in == 269) begin
					state<=10;
					out<=22;
				end
				if(in == 270) begin
					state<=10;
					out<=23;
				end
				if(in == 271) begin
					state<=10;
					out<=24;
				end
				if(in == 272) begin
					state<=10;
					out<=25;
				end
				if(in == 273) begin
					state<=10;
					out<=26;
				end
				if(in == 274) begin
					state<=10;
					out<=27;
				end
				if(in == 275) begin
					state<=10;
					out<=28;
				end
				if(in == 276) begin
					state<=10;
					out<=29;
				end
				if(in == 277) begin
					state<=10;
					out<=30;
				end
				if(in == 278) begin
					state<=10;
					out<=31;
				end
				if(in == 279) begin
					state<=10;
					out<=32;
				end
				if(in == 280) begin
					state<=10;
					out<=33;
				end
				if(in == 281) begin
					state<=10;
					out<=34;
				end
				if(in == 282) begin
					state<=10;
					out<=35;
				end
				if(in == 283) begin
					state<=10;
					out<=36;
				end
				if(in == 284) begin
					state<=10;
					out<=37;
				end
				if(in == 285) begin
					state<=3;
					out<=38;
				end
				if(in == 286) begin
					state<=9;
					out<=39;
				end
				if(in == 287) begin
					state<=3;
					out<=40;
				end
				if(in == 288) begin
					state<=10;
					out<=41;
				end
				if(in == 289) begin
					state<=3;
					out<=42;
				end
				if(in == 290) begin
					state<=10;
					out<=43;
				end
				if(in == 291) begin
					state<=10;
					out<=44;
				end
				if(in == 292) begin
					state<=10;
					out<=45;
				end
				if(in == 293) begin
					state<=10;
					out<=46;
				end
				if(in == 294) begin
					state<=10;
					out<=47;
				end
				if(in == 295) begin
					state<=10;
					out<=48;
				end
				if(in == 296) begin
					state<=10;
					out<=49;
				end
				if(in == 297) begin
					state<=10;
					out<=50;
				end
				if(in == 298) begin
					state<=10;
					out<=51;
				end
				if(in == 299) begin
					state<=10;
					out<=52;
				end
				if(in == 300) begin
					state<=10;
					out<=53;
				end
				if(in == 301) begin
					state<=10;
					out<=54;
				end
				if(in == 302) begin
					state<=10;
					out<=55;
				end
				if(in == 303) begin
					state<=10;
					out<=56;
				end
				if(in == 304) begin
					state<=10;
					out<=57;
				end
				if(in == 305) begin
					state<=10;
					out<=58;
				end
				if(in == 306) begin
					state<=10;
					out<=59;
				end
				if(in == 307) begin
					state<=10;
					out<=60;
				end
				if(in == 308) begin
					state<=10;
					out<=61;
				end
				if(in == 309) begin
					state<=10;
					out<=62;
				end
				if(in == 310) begin
					state<=10;
					out<=63;
				end
				if(in == 311) begin
					state<=10;
					out<=64;
				end
				if(in == 312) begin
					state<=10;
					out<=65;
				end
				if(in == 313) begin
					state<=10;
					out<=66;
				end
				if(in == 314) begin
					state<=10;
					out<=67;
				end
				if(in == 315) begin
					state<=10;
					out<=68;
				end
				if(in == 316) begin
					state<=10;
					out<=69;
				end
				if(in == 317) begin
					state<=10;
					out<=70;
				end
				if(in == 318) begin
					state<=10;
					out<=71;
				end
				if(in == 319) begin
					state<=10;
					out<=72;
				end
				if(in == 320) begin
					state<=10;
					out<=73;
				end
				if(in == 321) begin
					state<=10;
					out<=74;
				end
				if(in == 322) begin
					state<=10;
					out<=75;
				end
				if(in == 323) begin
					state<=10;
					out<=76;
				end
				if(in == 324) begin
					state<=10;
					out<=77;
				end
				if(in == 325) begin
					state<=10;
					out<=78;
				end
				if(in == 326) begin
					state<=10;
					out<=79;
				end
				if(in == 327) begin
					state<=10;
					out<=80;
				end
				if(in == 328) begin
					state<=10;
					out<=81;
				end
				if(in == 329) begin
					state<=10;
					out<=82;
				end
				if(in == 330) begin
					state<=10;
					out<=83;
				end
				if(in == 331) begin
					state<=10;
					out<=84;
				end
				if(in == 332) begin
					state<=10;
					out<=85;
				end
				if(in == 333) begin
					state<=10;
					out<=86;
				end
				if(in == 334) begin
					state<=10;
					out<=87;
				end
				if(in == 335) begin
					state<=10;
					out<=88;
				end
				if(in == 336) begin
					state<=10;
					out<=89;
				end
				if(in == 337) begin
					state<=2;
					out<=90;
				end
				if(in == 338) begin
					state<=2;
					out<=91;
				end
				if(in == 339) begin
					state<=2;
					out<=92;
				end
				if(in == 340) begin
					state<=2;
					out<=93;
				end
				if(in == 341) begin
					state<=2;
					out<=94;
				end
				if(in == 342) begin
					state<=2;
					out<=95;
				end
				if(in == 343) begin
					state<=2;
					out<=96;
				end
				if(in == 344) begin
					state<=2;
					out<=97;
				end
				if(in == 345) begin
					state<=2;
					out<=98;
				end
				if(in == 346) begin
					state<=2;
					out<=99;
				end
				if(in == 347) begin
					state<=2;
					out<=100;
				end
				if(in == 348) begin
					state<=2;
					out<=101;
				end
				if(in == 349) begin
					state<=3;
					out<=102;
				end
				if(in == 350) begin
					state<=9;
					out<=103;
				end
				if(in == 351) begin
					state<=3;
					out<=104;
				end
				if(in == 352) begin
					state<=10;
					out<=105;
				end
				if(in == 353) begin
					state<=3;
					out<=106;
				end
				if(in == 354) begin
					state<=10;
					out<=107;
				end
				if(in == 355) begin
					state<=10;
					out<=108;
				end
				if(in == 356) begin
					state<=10;
					out<=109;
				end
				if(in == 357) begin
					state<=10;
					out<=110;
				end
				if(in == 358) begin
					state<=10;
					out<=111;
				end
				if(in == 359) begin
					state<=10;
					out<=112;
				end
				if(in == 360) begin
					state<=10;
					out<=113;
				end
				if(in == 361) begin
					state<=10;
					out<=114;
				end
				if(in == 362) begin
					state<=10;
					out<=115;
				end
				if(in == 363) begin
					state<=10;
					out<=116;
				end
				if(in == 364) begin
					state<=10;
					out<=117;
				end
				if(in == 365) begin
					state<=10;
					out<=118;
				end
				if(in == 366) begin
					state<=10;
					out<=119;
				end
				if(in == 367) begin
					state<=10;
					out<=120;
				end
				if(in == 368) begin
					state<=10;
					out<=121;
				end
				if(in == 369) begin
					state<=10;
					out<=122;
				end
				if(in == 370) begin
					state<=10;
					out<=123;
				end
				if(in == 371) begin
					state<=10;
					out<=124;
				end
				if(in == 372) begin
					state<=10;
					out<=125;
				end
				if(in == 373) begin
					state<=10;
					out<=126;
				end
				if(in == 374) begin
					state<=10;
					out<=127;
				end
				if(in == 375) begin
					state<=10;
					out<=128;
				end
				if(in == 376) begin
					state<=10;
					out<=129;
				end
				if(in == 377) begin
					state<=10;
					out<=130;
				end
				if(in == 378) begin
					state<=10;
					out<=131;
				end
				if(in == 379) begin
					state<=10;
					out<=132;
				end
				if(in == 380) begin
					state<=10;
					out<=133;
				end
				if(in == 381) begin
					state<=10;
					out<=134;
				end
				if(in == 382) begin
					state<=10;
					out<=135;
				end
				if(in == 383) begin
					state<=10;
					out<=136;
				end
				if(in == 384) begin
					state<=10;
					out<=137;
				end
				if(in == 385) begin
					state<=10;
					out<=138;
				end
				if(in == 386) begin
					state<=10;
					out<=139;
				end
				if(in == 387) begin
					state<=10;
					out<=140;
				end
				if(in == 388) begin
					state<=10;
					out<=141;
				end
				if(in == 389) begin
					state<=10;
					out<=142;
				end
				if(in == 390) begin
					state<=10;
					out<=143;
				end
				if(in == 391) begin
					state<=10;
					out<=144;
				end
				if(in == 392) begin
					state<=10;
					out<=145;
				end
				if(in == 393) begin
					state<=10;
					out<=146;
				end
				if(in == 394) begin
					state<=10;
					out<=147;
				end
				if(in == 395) begin
					state<=10;
					out<=148;
				end
				if(in == 396) begin
					state<=10;
					out<=149;
				end
				if(in == 397) begin
					state<=10;
					out<=150;
				end
				if(in == 398) begin
					state<=10;
					out<=151;
				end
				if(in == 399) begin
					state<=10;
					out<=152;
				end
				if(in == 400) begin
					state<=10;
					out<=153;
				end
				if(in == 401) begin
					state<=3;
					out<=154;
				end
				if(in == 402) begin
					state<=9;
					out<=155;
				end
				if(in == 403) begin
					state<=3;
					out<=156;
				end
				if(in == 404) begin
					state<=10;
					out<=157;
				end
				if(in == 405) begin
					state<=3;
					out<=158;
				end
				if(in == 406) begin
					state<=10;
					out<=159;
				end
				if(in == 407) begin
					state<=10;
					out<=160;
				end
				if(in == 408) begin
					state<=10;
					out<=161;
				end
				if(in == 409) begin
					state<=10;
					out<=162;
				end
				if(in == 410) begin
					state<=10;
					out<=163;
				end
				if(in == 411) begin
					state<=10;
					out<=164;
				end
				if(in == 412) begin
					state<=10;
					out<=165;
				end
				if(in == 413) begin
					state<=10;
					out<=166;
				end
				if(in == 414) begin
					state<=10;
					out<=167;
				end
				if(in == 415) begin
					state<=10;
					out<=168;
				end
				if(in == 416) begin
					state<=10;
					out<=169;
				end
				if(in == 417) begin
					state<=10;
					out<=170;
				end
				if(in == 418) begin
					state<=10;
					out<=171;
				end
				if(in == 419) begin
					state<=10;
					out<=172;
				end
				if(in == 420) begin
					state<=10;
					out<=173;
				end
				if(in == 421) begin
					state<=10;
					out<=174;
				end
				if(in == 422) begin
					state<=10;
					out<=175;
				end
				if(in == 423) begin
					state<=10;
					out<=176;
				end
				if(in == 424) begin
					state<=10;
					out<=177;
				end
				if(in == 425) begin
					state<=10;
					out<=178;
				end
				if(in == 426) begin
					state<=10;
					out<=179;
				end
				if(in == 427) begin
					state<=10;
					out<=180;
				end
				if(in == 428) begin
					state<=10;
					out<=181;
				end
				if(in == 429) begin
					state<=10;
					out<=182;
				end
				if(in == 430) begin
					state<=10;
					out<=183;
				end
				if(in == 431) begin
					state<=10;
					out<=184;
				end
				if(in == 432) begin
					state<=10;
					out<=185;
				end
				if(in == 433) begin
					state<=10;
					out<=186;
				end
				if(in == 434) begin
					state<=10;
					out<=187;
				end
				if(in == 435) begin
					state<=10;
					out<=188;
				end
				if(in == 436) begin
					state<=10;
					out<=189;
				end
				if(in == 437) begin
					state<=10;
					out<=190;
				end
				if(in == 438) begin
					state<=10;
					out<=191;
				end
				if(in == 439) begin
					state<=10;
					out<=192;
				end
				if(in == 440) begin
					state<=10;
					out<=193;
				end
				if(in == 441) begin
					state<=10;
					out<=194;
				end
				if(in == 442) begin
					state<=10;
					out<=195;
				end
				if(in == 443) begin
					state<=10;
					out<=196;
				end
				if(in == 444) begin
					state<=10;
					out<=197;
				end
				if(in == 445) begin
					state<=10;
					out<=198;
				end
				if(in == 446) begin
					state<=10;
					out<=199;
				end
				if(in == 447) begin
					state<=10;
					out<=200;
				end
				if(in == 448) begin
					state<=10;
					out<=201;
				end
				if(in == 449) begin
					state<=10;
					out<=202;
				end
				if(in == 450) begin
					state<=10;
					out<=203;
				end
				if(in == 451) begin
					state<=10;
					out<=204;
				end
				if(in == 452) begin
					state<=10;
					out<=205;
				end
				if(in == 453) begin
					state<=2;
					out<=206;
				end
				if(in == 454) begin
					state<=2;
					out<=207;
				end
				if(in == 455) begin
					state<=2;
					out<=208;
				end
				if(in == 456) begin
					state<=2;
					out<=209;
				end
				if(in == 457) begin
					state<=2;
					out<=210;
				end
				if(in == 458) begin
					state<=2;
					out<=211;
				end
				if(in == 459) begin
					state<=2;
					out<=212;
				end
				if(in == 460) begin
					state<=2;
					out<=213;
				end
				if(in == 461) begin
					state<=2;
					out<=214;
				end
				if(in == 462) begin
					state<=2;
					out<=215;
				end
				if(in == 463) begin
					state<=2;
					out<=216;
				end
				if(in == 464) begin
					state<=2;
					out<=217;
				end
				if(in == 465) begin
					state<=3;
					out<=218;
				end
				if(in == 466) begin
					state<=9;
					out<=219;
				end
				if(in == 467) begin
					state<=3;
					out<=220;
				end
				if(in == 468) begin
					state<=10;
					out<=221;
				end
				if(in == 469) begin
					state<=3;
					out<=222;
				end
				if(in == 470) begin
					state<=10;
					out<=223;
				end
				if(in == 471) begin
					state<=10;
					out<=224;
				end
				if(in == 472) begin
					state<=10;
					out<=225;
				end
				if(in == 473) begin
					state<=10;
					out<=226;
				end
				if(in == 474) begin
					state<=10;
					out<=227;
				end
				if(in == 475) begin
					state<=10;
					out<=228;
				end
				if(in == 476) begin
					state<=10;
					out<=229;
				end
				if(in == 477) begin
					state<=10;
					out<=230;
				end
				if(in == 478) begin
					state<=10;
					out<=231;
				end
				if(in == 479) begin
					state<=10;
					out<=232;
				end
				if(in == 480) begin
					state<=10;
					out<=233;
				end
				if(in == 481) begin
					state<=10;
					out<=234;
				end
				if(in == 482) begin
					state<=10;
					out<=235;
				end
				if(in == 483) begin
					state<=10;
					out<=236;
				end
				if(in == 484) begin
					state<=10;
					out<=237;
				end
				if(in == 485) begin
					state<=10;
					out<=238;
				end
				if(in == 486) begin
					state<=10;
					out<=239;
				end
				if(in == 487) begin
					state<=10;
					out<=240;
				end
				if(in == 488) begin
					state<=10;
					out<=241;
				end
				if(in == 489) begin
					state<=10;
					out<=242;
				end
				if(in == 490) begin
					state<=10;
					out<=243;
				end
				if(in == 491) begin
					state<=10;
					out<=244;
				end
				if(in == 492) begin
					state<=10;
					out<=245;
				end
				if(in == 493) begin
					state<=10;
					out<=246;
				end
				if(in == 494) begin
					state<=10;
					out<=247;
				end
				if(in == 495) begin
					state<=10;
					out<=248;
				end
				if(in == 496) begin
					state<=10;
					out<=249;
				end
				if(in == 497) begin
					state<=10;
					out<=250;
				end
				if(in == 498) begin
					state<=10;
					out<=251;
				end
				if(in == 499) begin
					state<=10;
					out<=252;
				end
				if(in == 500) begin
					state<=10;
					out<=253;
				end
				if(in == 501) begin
					state<=10;
					out<=254;
				end
				if(in == 502) begin
					state<=10;
					out<=255;
				end
				if(in == 503) begin
					state<=10;
					out<=0;
				end
				if(in == 504) begin
					state<=10;
					out<=1;
				end
				if(in == 505) begin
					state<=10;
					out<=2;
				end
				if(in == 506) begin
					state<=10;
					out<=3;
				end
				if(in == 507) begin
					state<=10;
					out<=4;
				end
				if(in == 508) begin
					state<=10;
					out<=5;
				end
				if(in == 509) begin
					state<=10;
					out<=6;
				end
				if(in == 510) begin
					state<=10;
					out<=7;
				end
				if(in == 511) begin
					state<=10;
					out<=8;
				end
				if(in == 512) begin
					state<=10;
					out<=9;
				end
				if(in == 513) begin
					state<=10;
					out<=10;
				end
				if(in == 514) begin
					state<=10;
					out<=11;
				end
				if(in == 515) begin
					state<=10;
					out<=12;
				end
				if(in == 516) begin
					state<=10;
					out<=13;
				end
				if(in == 517) begin
					state<=3;
					out<=14;
				end
				if(in == 518) begin
					state<=9;
					out<=15;
				end
				if(in == 519) begin
					state<=3;
					out<=16;
				end
				if(in == 520) begin
					state<=10;
					out<=17;
				end
				if(in == 521) begin
					state<=3;
					out<=18;
				end
				if(in == 522) begin
					state<=10;
					out<=19;
				end
				if(in == 523) begin
					state<=10;
					out<=20;
				end
				if(in == 524) begin
					state<=10;
					out<=21;
				end
				if(in == 525) begin
					state<=10;
					out<=22;
				end
				if(in == 526) begin
					state<=10;
					out<=23;
				end
				if(in == 527) begin
					state<=10;
					out<=24;
				end
				if(in == 528) begin
					state<=10;
					out<=25;
				end
				if(in == 529) begin
					state<=10;
					out<=26;
				end
				if(in == 530) begin
					state<=10;
					out<=27;
				end
				if(in == 531) begin
					state<=10;
					out<=28;
				end
				if(in == 532) begin
					state<=10;
					out<=29;
				end
				if(in == 533) begin
					state<=10;
					out<=30;
				end
				if(in == 534) begin
					state<=10;
					out<=31;
				end
				if(in == 535) begin
					state<=10;
					out<=32;
				end
				if(in == 536) begin
					state<=10;
					out<=33;
				end
				if(in == 537) begin
					state<=10;
					out<=34;
				end
				if(in == 538) begin
					state<=10;
					out<=35;
				end
				if(in == 539) begin
					state<=10;
					out<=36;
				end
				if(in == 540) begin
					state<=10;
					out<=37;
				end
				if(in == 541) begin
					state<=10;
					out<=38;
				end
				if(in == 542) begin
					state<=10;
					out<=39;
				end
				if(in == 543) begin
					state<=10;
					out<=40;
				end
				if(in == 544) begin
					state<=10;
					out<=41;
				end
				if(in == 545) begin
					state<=10;
					out<=42;
				end
				if(in == 546) begin
					state<=10;
					out<=43;
				end
				if(in == 547) begin
					state<=10;
					out<=44;
				end
				if(in == 548) begin
					state<=10;
					out<=45;
				end
				if(in == 549) begin
					state<=10;
					out<=46;
				end
				if(in == 550) begin
					state<=10;
					out<=47;
				end
				if(in == 551) begin
					state<=10;
					out<=48;
				end
				if(in == 552) begin
					state<=10;
					out<=49;
				end
				if(in == 553) begin
					state<=10;
					out<=50;
				end
				if(in == 554) begin
					state<=10;
					out<=51;
				end
				if(in == 555) begin
					state<=10;
					out<=52;
				end
				if(in == 556) begin
					state<=10;
					out<=53;
				end
				if(in == 557) begin
					state<=10;
					out<=54;
				end
				if(in == 558) begin
					state<=10;
					out<=55;
				end
				if(in == 559) begin
					state<=10;
					out<=56;
				end
				if(in == 560) begin
					state<=10;
					out<=57;
				end
				if(in == 561) begin
					state<=10;
					out<=58;
				end
				if(in == 562) begin
					state<=10;
					out<=59;
				end
				if(in == 563) begin
					state<=10;
					out<=60;
				end
				if(in == 564) begin
					state<=10;
					out<=61;
				end
				if(in == 565) begin
					state<=10;
					out<=62;
				end
				if(in == 566) begin
					state<=10;
					out<=63;
				end
				if(in == 567) begin
					state<=10;
					out<=64;
				end
				if(in == 568) begin
					state<=10;
					out<=65;
				end
				if(in == 569) begin
					state<=2;
					out<=66;
				end
				if(in == 570) begin
					state<=2;
					out<=67;
				end
				if(in == 571) begin
					state<=2;
					out<=68;
				end
				if(in == 572) begin
					state<=2;
					out<=69;
				end
				if(in == 573) begin
					state<=2;
					out<=70;
				end
				if(in == 574) begin
					state<=2;
					out<=71;
				end
				if(in == 575) begin
					state<=2;
					out<=72;
				end
				if(in == 576) begin
					state<=2;
					out<=73;
				end
				if(in == 577) begin
					state<=2;
					out<=74;
				end
				if(in == 578) begin
					state<=2;
					out<=75;
				end
				if(in == 579) begin
					state<=2;
					out<=76;
				end
				if(in == 580) begin
					state<=2;
					out<=77;
				end
				if(in == 581) begin
					state<=3;
					out<=78;
				end
				if(in == 582) begin
					state<=9;
					out<=79;
				end
				if(in == 583) begin
					state<=3;
					out<=80;
				end
				if(in == 584) begin
					state<=10;
					out<=81;
				end
				if(in == 585) begin
					state<=3;
					out<=82;
				end
				if(in == 586) begin
					state<=10;
					out<=83;
				end
				if(in == 587) begin
					state<=10;
					out<=84;
				end
				if(in == 588) begin
					state<=10;
					out<=85;
				end
				if(in == 589) begin
					state<=10;
					out<=86;
				end
				if(in == 590) begin
					state<=10;
					out<=87;
				end
				if(in == 591) begin
					state<=10;
					out<=88;
				end
				if(in == 592) begin
					state<=10;
					out<=89;
				end
				if(in == 593) begin
					state<=10;
					out<=90;
				end
				if(in == 594) begin
					state<=10;
					out<=91;
				end
				if(in == 595) begin
					state<=10;
					out<=92;
				end
				if(in == 596) begin
					state<=10;
					out<=93;
				end
				if(in == 597) begin
					state<=10;
					out<=94;
				end
				if(in == 598) begin
					state<=10;
					out<=95;
				end
				if(in == 599) begin
					state<=10;
					out<=96;
				end
				if(in == 600) begin
					state<=10;
					out<=97;
				end
				if(in == 601) begin
					state<=10;
					out<=98;
				end
				if(in == 602) begin
					state<=10;
					out<=99;
				end
				if(in == 603) begin
					state<=10;
					out<=100;
				end
				if(in == 604) begin
					state<=10;
					out<=101;
				end
				if(in == 605) begin
					state<=10;
					out<=102;
				end
				if(in == 606) begin
					state<=10;
					out<=103;
				end
				if(in == 607) begin
					state<=10;
					out<=104;
				end
				if(in == 608) begin
					state<=10;
					out<=105;
				end
				if(in == 609) begin
					state<=10;
					out<=106;
				end
				if(in == 610) begin
					state<=10;
					out<=107;
				end
				if(in == 611) begin
					state<=10;
					out<=108;
				end
				if(in == 612) begin
					state<=10;
					out<=109;
				end
				if(in == 613) begin
					state<=10;
					out<=110;
				end
				if(in == 614) begin
					state<=10;
					out<=111;
				end
				if(in == 615) begin
					state<=10;
					out<=112;
				end
				if(in == 616) begin
					state<=10;
					out<=113;
				end
				if(in == 617) begin
					state<=10;
					out<=114;
				end
				if(in == 618) begin
					state<=10;
					out<=115;
				end
				if(in == 619) begin
					state<=10;
					out<=116;
				end
				if(in == 620) begin
					state<=10;
					out<=117;
				end
				if(in == 621) begin
					state<=10;
					out<=118;
				end
				if(in == 622) begin
					state<=10;
					out<=119;
				end
				if(in == 623) begin
					state<=10;
					out<=120;
				end
				if(in == 624) begin
					state<=10;
					out<=121;
				end
				if(in == 625) begin
					state<=10;
					out<=122;
				end
				if(in == 626) begin
					state<=10;
					out<=123;
				end
				if(in == 627) begin
					state<=10;
					out<=124;
				end
				if(in == 628) begin
					state<=10;
					out<=125;
				end
				if(in == 629) begin
					state<=10;
					out<=126;
				end
				if(in == 630) begin
					state<=10;
					out<=127;
				end
				if(in == 631) begin
					state<=10;
					out<=128;
				end
				if(in == 632) begin
					state<=10;
					out<=129;
				end
				if(in == 633) begin
					state<=3;
					out<=130;
				end
				if(in == 634) begin
					state<=9;
					out<=131;
				end
				if(in == 635) begin
					state<=3;
					out<=132;
				end
				if(in == 636) begin
					state<=10;
					out<=133;
				end
				if(in == 637) begin
					state<=3;
					out<=134;
				end
				if(in == 638) begin
					state<=10;
					out<=135;
				end
				if(in == 639) begin
					state<=10;
					out<=136;
				end
				if(in == 640) begin
					state<=10;
					out<=137;
				end
				if(in == 641) begin
					state<=10;
					out<=138;
				end
				if(in == 642) begin
					state<=10;
					out<=139;
				end
				if(in == 643) begin
					state<=10;
					out<=140;
				end
				if(in == 644) begin
					state<=10;
					out<=141;
				end
				if(in == 645) begin
					state<=10;
					out<=142;
				end
				if(in == 646) begin
					state<=10;
					out<=143;
				end
				if(in == 647) begin
					state<=10;
					out<=144;
				end
				if(in == 648) begin
					state<=10;
					out<=145;
				end
				if(in == 649) begin
					state<=10;
					out<=146;
				end
				if(in == 650) begin
					state<=10;
					out<=147;
				end
				if(in == 651) begin
					state<=10;
					out<=148;
				end
				if(in == 652) begin
					state<=10;
					out<=149;
				end
				if(in == 653) begin
					state<=10;
					out<=150;
				end
				if(in == 654) begin
					state<=10;
					out<=151;
				end
				if(in == 655) begin
					state<=10;
					out<=152;
				end
				if(in == 656) begin
					state<=10;
					out<=153;
				end
				if(in == 657) begin
					state<=10;
					out<=154;
				end
				if(in == 658) begin
					state<=10;
					out<=155;
				end
				if(in == 659) begin
					state<=10;
					out<=156;
				end
				if(in == 660) begin
					state<=10;
					out<=157;
				end
				if(in == 661) begin
					state<=10;
					out<=158;
				end
				if(in == 662) begin
					state<=10;
					out<=159;
				end
				if(in == 663) begin
					state<=10;
					out<=160;
				end
				if(in == 664) begin
					state<=10;
					out<=161;
				end
				if(in == 665) begin
					state<=10;
					out<=162;
				end
				if(in == 666) begin
					state<=10;
					out<=163;
				end
				if(in == 667) begin
					state<=10;
					out<=164;
				end
				if(in == 668) begin
					state<=10;
					out<=165;
				end
				if(in == 669) begin
					state<=10;
					out<=166;
				end
				if(in == 670) begin
					state<=10;
					out<=167;
				end
				if(in == 671) begin
					state<=10;
					out<=168;
				end
				if(in == 672) begin
					state<=10;
					out<=169;
				end
				if(in == 673) begin
					state<=10;
					out<=170;
				end
				if(in == 674) begin
					state<=10;
					out<=171;
				end
				if(in == 675) begin
					state<=10;
					out<=172;
				end
				if(in == 676) begin
					state<=10;
					out<=173;
				end
				if(in == 677) begin
					state<=10;
					out<=174;
				end
				if(in == 678) begin
					state<=10;
					out<=175;
				end
				if(in == 679) begin
					state<=10;
					out<=176;
				end
				if(in == 680) begin
					state<=10;
					out<=177;
				end
				if(in == 681) begin
					state<=10;
					out<=178;
				end
				if(in == 682) begin
					state<=10;
					out<=179;
				end
				if(in == 683) begin
					state<=10;
					out<=180;
				end
				if(in == 684) begin
					state<=10;
					out<=181;
				end
				if(in == 685) begin
					state<=2;
					out<=182;
				end
				if(in == 686) begin
					state<=2;
					out<=183;
				end
				if(in == 687) begin
					state<=2;
					out<=184;
				end
				if(in == 688) begin
					state<=2;
					out<=185;
				end
				if(in == 689) begin
					state<=2;
					out<=186;
				end
				if(in == 690) begin
					state<=2;
					out<=187;
				end
				if(in == 691) begin
					state<=2;
					out<=188;
				end
				if(in == 692) begin
					state<=2;
					out<=189;
				end
				if(in == 693) begin
					state<=2;
					out<=190;
				end
				if(in == 694) begin
					state<=2;
					out<=191;
				end
				if(in == 695) begin
					state<=2;
					out<=192;
				end
				if(in == 696) begin
					state<=2;
					out<=193;
				end
				if(in == 697) begin
					state<=3;
					out<=194;
				end
				if(in == 698) begin
					state<=9;
					out<=195;
				end
				if(in == 699) begin
					state<=3;
					out<=196;
				end
				if(in == 700) begin
					state<=10;
					out<=197;
				end
				if(in == 701) begin
					state<=3;
					out<=198;
				end
				if(in == 702) begin
					state<=10;
					out<=199;
				end
				if(in == 703) begin
					state<=10;
					out<=200;
				end
				if(in == 704) begin
					state<=10;
					out<=201;
				end
				if(in == 705) begin
					state<=10;
					out<=202;
				end
				if(in == 706) begin
					state<=10;
					out<=203;
				end
				if(in == 707) begin
					state<=10;
					out<=204;
				end
				if(in == 708) begin
					state<=10;
					out<=205;
				end
				if(in == 709) begin
					state<=10;
					out<=206;
				end
				if(in == 710) begin
					state<=10;
					out<=207;
				end
				if(in == 711) begin
					state<=10;
					out<=208;
				end
				if(in == 712) begin
					state<=10;
					out<=209;
				end
				if(in == 713) begin
					state<=10;
					out<=210;
				end
				if(in == 714) begin
					state<=10;
					out<=211;
				end
				if(in == 715) begin
					state<=10;
					out<=212;
				end
				if(in == 716) begin
					state<=10;
					out<=213;
				end
				if(in == 717) begin
					state<=10;
					out<=214;
				end
				if(in == 718) begin
					state<=10;
					out<=215;
				end
				if(in == 719) begin
					state<=10;
					out<=216;
				end
				if(in == 720) begin
					state<=10;
					out<=217;
				end
				if(in == 721) begin
					state<=10;
					out<=218;
				end
				if(in == 722) begin
					state<=10;
					out<=219;
				end
				if(in == 723) begin
					state<=10;
					out<=220;
				end
				if(in == 724) begin
					state<=10;
					out<=221;
				end
				if(in == 725) begin
					state<=10;
					out<=222;
				end
				if(in == 726) begin
					state<=10;
					out<=223;
				end
				if(in == 727) begin
					state<=10;
					out<=224;
				end
				if(in == 728) begin
					state<=10;
					out<=225;
				end
				if(in == 729) begin
					state<=10;
					out<=226;
				end
				if(in == 730) begin
					state<=10;
					out<=227;
				end
				if(in == 731) begin
					state<=10;
					out<=228;
				end
				if(in == 732) begin
					state<=10;
					out<=229;
				end
				if(in == 733) begin
					state<=10;
					out<=230;
				end
				if(in == 734) begin
					state<=10;
					out<=231;
				end
				if(in == 735) begin
					state<=10;
					out<=232;
				end
				if(in == 736) begin
					state<=10;
					out<=233;
				end
				if(in == 737) begin
					state<=10;
					out<=234;
				end
				if(in == 738) begin
					state<=10;
					out<=235;
				end
				if(in == 739) begin
					state<=10;
					out<=236;
				end
				if(in == 740) begin
					state<=10;
					out<=237;
				end
				if(in == 741) begin
					state<=10;
					out<=238;
				end
				if(in == 742) begin
					state<=10;
					out<=239;
				end
				if(in == 743) begin
					state<=10;
					out<=240;
				end
				if(in == 744) begin
					state<=10;
					out<=241;
				end
				if(in == 745) begin
					state<=10;
					out<=242;
				end
				if(in == 746) begin
					state<=10;
					out<=243;
				end
				if(in == 747) begin
					state<=10;
					out<=244;
				end
				if(in == 748) begin
					state<=10;
					out<=245;
				end
				if(in == 749) begin
					state<=3;
					out<=246;
				end
				if(in == 750) begin
					state<=9;
					out<=247;
				end
				if(in == 751) begin
					state<=3;
					out<=248;
				end
				if(in == 752) begin
					state<=10;
					out<=249;
				end
				if(in == 753) begin
					state<=3;
					out<=250;
				end
				if(in == 754) begin
					state<=10;
					out<=251;
				end
				if(in == 755) begin
					state<=10;
					out<=252;
				end
				if(in == 756) begin
					state<=10;
					out<=253;
				end
				if(in == 757) begin
					state<=10;
					out<=254;
				end
				if(in == 758) begin
					state<=10;
					out<=255;
				end
				if(in == 759) begin
					state<=10;
					out<=0;
				end
				if(in == 760) begin
					state<=10;
					out<=1;
				end
				if(in == 761) begin
					state<=10;
					out<=2;
				end
				if(in == 762) begin
					state<=10;
					out<=3;
				end
				if(in == 763) begin
					state<=10;
					out<=4;
				end
				if(in == 764) begin
					state<=10;
					out<=5;
				end
				if(in == 765) begin
					state<=10;
					out<=6;
				end
				if(in == 766) begin
					state<=10;
					out<=7;
				end
				if(in == 767) begin
					state<=10;
					out<=8;
				end
				if(in == 768) begin
					state<=10;
					out<=9;
				end
				if(in == 769) begin
					state<=10;
					out<=10;
				end
				if(in == 770) begin
					state<=10;
					out<=11;
				end
				if(in == 771) begin
					state<=10;
					out<=12;
				end
				if(in == 772) begin
					state<=10;
					out<=13;
				end
				if(in == 773) begin
					state<=10;
					out<=14;
				end
				if(in == 774) begin
					state<=10;
					out<=15;
				end
				if(in == 775) begin
					state<=10;
					out<=16;
				end
				if(in == 776) begin
					state<=10;
					out<=17;
				end
				if(in == 777) begin
					state<=10;
					out<=18;
				end
				if(in == 778) begin
					state<=10;
					out<=19;
				end
				if(in == 779) begin
					state<=10;
					out<=20;
				end
				if(in == 780) begin
					state<=10;
					out<=21;
				end
				if(in == 781) begin
					state<=10;
					out<=22;
				end
				if(in == 782) begin
					state<=10;
					out<=23;
				end
				if(in == 783) begin
					state<=10;
					out<=24;
				end
				if(in == 784) begin
					state<=10;
					out<=25;
				end
				if(in == 785) begin
					state<=10;
					out<=26;
				end
				if(in == 786) begin
					state<=10;
					out<=27;
				end
				if(in == 787) begin
					state<=10;
					out<=28;
				end
				if(in == 788) begin
					state<=10;
					out<=29;
				end
				if(in == 789) begin
					state<=10;
					out<=30;
				end
				if(in == 790) begin
					state<=10;
					out<=31;
				end
				if(in == 791) begin
					state<=10;
					out<=32;
				end
				if(in == 792) begin
					state<=10;
					out<=33;
				end
				if(in == 793) begin
					state<=10;
					out<=34;
				end
				if(in == 794) begin
					state<=10;
					out<=35;
				end
				if(in == 795) begin
					state<=10;
					out<=36;
				end
				if(in == 796) begin
					state<=10;
					out<=37;
				end
				if(in == 797) begin
					state<=10;
					out<=38;
				end
				if(in == 798) begin
					state<=10;
					out<=39;
				end
				if(in == 799) begin
					state<=10;
					out<=40;
				end
				if(in == 800) begin
					state<=10;
					out<=41;
				end
				if(in == 801) begin
					state<=2;
					out<=42;
				end
				if(in == 802) begin
					state<=2;
					out<=43;
				end
				if(in == 803) begin
					state<=2;
					out<=44;
				end
				if(in == 804) begin
					state<=2;
					out<=45;
				end
				if(in == 805) begin
					state<=2;
					out<=46;
				end
				if(in == 806) begin
					state<=2;
					out<=47;
				end
				if(in == 807) begin
					state<=2;
					out<=48;
				end
				if(in == 808) begin
					state<=2;
					out<=49;
				end
				if(in == 809) begin
					state<=2;
					out<=50;
				end
				if(in == 810) begin
					state<=2;
					out<=51;
				end
				if(in == 811) begin
					state<=2;
					out<=52;
				end
				if(in == 812) begin
					state<=2;
					out<=53;
				end
				if(in == 813) begin
					state<=3;
					out<=54;
				end
				if(in == 814) begin
					state<=9;
					out<=55;
				end
				if(in == 815) begin
					state<=3;
					out<=56;
				end
				if(in == 816) begin
					state<=10;
					out<=57;
				end
				if(in == 817) begin
					state<=3;
					out<=58;
				end
				if(in == 818) begin
					state<=10;
					out<=59;
				end
				if(in == 819) begin
					state<=10;
					out<=60;
				end
				if(in == 820) begin
					state<=10;
					out<=61;
				end
				if(in == 821) begin
					state<=10;
					out<=62;
				end
				if(in == 822) begin
					state<=10;
					out<=63;
				end
				if(in == 823) begin
					state<=10;
					out<=64;
				end
				if(in == 824) begin
					state<=10;
					out<=65;
				end
				if(in == 825) begin
					state<=10;
					out<=66;
				end
				if(in == 826) begin
					state<=10;
					out<=67;
				end
				if(in == 827) begin
					state<=10;
					out<=68;
				end
				if(in == 828) begin
					state<=10;
					out<=69;
				end
				if(in == 829) begin
					state<=10;
					out<=70;
				end
				if(in == 830) begin
					state<=10;
					out<=71;
				end
				if(in == 831) begin
					state<=10;
					out<=72;
				end
				if(in == 832) begin
					state<=10;
					out<=73;
				end
				if(in == 833) begin
					state<=10;
					out<=74;
				end
				if(in == 834) begin
					state<=10;
					out<=75;
				end
				if(in == 835) begin
					state<=10;
					out<=76;
				end
				if(in == 836) begin
					state<=10;
					out<=77;
				end
				if(in == 837) begin
					state<=10;
					out<=78;
				end
				if(in == 838) begin
					state<=10;
					out<=79;
				end
				if(in == 839) begin
					state<=10;
					out<=80;
				end
				if(in == 840) begin
					state<=10;
					out<=81;
				end
				if(in == 841) begin
					state<=10;
					out<=82;
				end
				if(in == 842) begin
					state<=10;
					out<=83;
				end
				if(in == 843) begin
					state<=10;
					out<=84;
				end
				if(in == 844) begin
					state<=10;
					out<=85;
				end
				if(in == 845) begin
					state<=10;
					out<=86;
				end
				if(in == 846) begin
					state<=10;
					out<=87;
				end
				if(in == 847) begin
					state<=10;
					out<=88;
				end
				if(in == 848) begin
					state<=10;
					out<=89;
				end
				if(in == 849) begin
					state<=10;
					out<=90;
				end
				if(in == 850) begin
					state<=10;
					out<=91;
				end
				if(in == 851) begin
					state<=10;
					out<=92;
				end
				if(in == 852) begin
					state<=10;
					out<=93;
				end
				if(in == 853) begin
					state<=10;
					out<=94;
				end
				if(in == 854) begin
					state<=10;
					out<=95;
				end
				if(in == 855) begin
					state<=10;
					out<=96;
				end
				if(in == 856) begin
					state<=10;
					out<=97;
				end
				if(in == 857) begin
					state<=10;
					out<=98;
				end
				if(in == 858) begin
					state<=10;
					out<=99;
				end
				if(in == 859) begin
					state<=10;
					out<=100;
				end
				if(in == 860) begin
					state<=10;
					out<=101;
				end
				if(in == 861) begin
					state<=10;
					out<=102;
				end
				if(in == 862) begin
					state<=10;
					out<=103;
				end
				if(in == 863) begin
					state<=10;
					out<=104;
				end
				if(in == 864) begin
					state<=10;
					out<=105;
				end
				if(in == 865) begin
					state<=3;
					out<=106;
				end
				if(in == 866) begin
					state<=9;
					out<=107;
				end
				if(in == 867) begin
					state<=3;
					out<=108;
				end
				if(in == 868) begin
					state<=10;
					out<=109;
				end
				if(in == 869) begin
					state<=3;
					out<=110;
				end
				if(in == 870) begin
					state<=10;
					out<=111;
				end
				if(in == 871) begin
					state<=10;
					out<=112;
				end
				if(in == 872) begin
					state<=10;
					out<=113;
				end
				if(in == 873) begin
					state<=10;
					out<=114;
				end
				if(in == 874) begin
					state<=10;
					out<=115;
				end
				if(in == 875) begin
					state<=10;
					out<=116;
				end
				if(in == 876) begin
					state<=10;
					out<=117;
				end
				if(in == 877) begin
					state<=10;
					out<=118;
				end
				if(in == 878) begin
					state<=10;
					out<=119;
				end
				if(in == 879) begin
					state<=10;
					out<=120;
				end
				if(in == 880) begin
					state<=10;
					out<=121;
				end
				if(in == 881) begin
					state<=10;
					out<=122;
				end
				if(in == 882) begin
					state<=10;
					out<=123;
				end
				if(in == 883) begin
					state<=10;
					out<=124;
				end
				if(in == 884) begin
					state<=10;
					out<=125;
				end
				if(in == 885) begin
					state<=10;
					out<=126;
				end
				if(in == 886) begin
					state<=10;
					out<=127;
				end
				if(in == 887) begin
					state<=10;
					out<=128;
				end
				if(in == 888) begin
					state<=10;
					out<=129;
				end
				if(in == 889) begin
					state<=10;
					out<=130;
				end
				if(in == 890) begin
					state<=10;
					out<=131;
				end
				if(in == 891) begin
					state<=10;
					out<=132;
				end
				if(in == 892) begin
					state<=10;
					out<=133;
				end
				if(in == 893) begin
					state<=10;
					out<=134;
				end
				if(in == 894) begin
					state<=10;
					out<=135;
				end
				if(in == 895) begin
					state<=10;
					out<=136;
				end
				if(in == 896) begin
					state<=10;
					out<=137;
				end
				if(in == 897) begin
					state<=10;
					out<=138;
				end
				if(in == 898) begin
					state<=10;
					out<=139;
				end
				if(in == 899) begin
					state<=10;
					out<=140;
				end
				if(in == 900) begin
					state<=10;
					out<=141;
				end
				if(in == 901) begin
					state<=10;
					out<=142;
				end
				if(in == 902) begin
					state<=10;
					out<=143;
				end
				if(in == 903) begin
					state<=10;
					out<=144;
				end
				if(in == 904) begin
					state<=10;
					out<=145;
				end
				if(in == 905) begin
					state<=10;
					out<=146;
				end
				if(in == 906) begin
					state<=10;
					out<=147;
				end
				if(in == 907) begin
					state<=10;
					out<=148;
				end
				if(in == 908) begin
					state<=10;
					out<=149;
				end
				if(in == 909) begin
					state<=10;
					out<=150;
				end
				if(in == 910) begin
					state<=10;
					out<=151;
				end
				if(in == 911) begin
					state<=10;
					out<=152;
				end
				if(in == 912) begin
					state<=10;
					out<=153;
				end
				if(in == 913) begin
					state<=10;
					out<=154;
				end
				if(in == 914) begin
					state<=10;
					out<=155;
				end
				if(in == 915) begin
					state<=10;
					out<=156;
				end
				if(in == 916) begin
					state<=10;
					out<=157;
				end
				if(in == 917) begin
					state<=2;
					out<=158;
				end
				if(in == 918) begin
					state<=2;
					out<=159;
				end
				if(in == 919) begin
					state<=2;
					out<=160;
				end
				if(in == 920) begin
					state<=2;
					out<=161;
				end
				if(in == 921) begin
					state<=2;
					out<=162;
				end
				if(in == 922) begin
					state<=2;
					out<=163;
				end
				if(in == 923) begin
					state<=2;
					out<=164;
				end
				if(in == 924) begin
					state<=2;
					out<=165;
				end
				if(in == 925) begin
					state<=2;
					out<=166;
				end
				if(in == 926) begin
					state<=2;
					out<=167;
				end
				if(in == 927) begin
					state<=2;
					out<=168;
				end
				if(in == 928) begin
					state<=2;
					out<=169;
				end
			end
			10: begin
				if(in == 0) begin
					state<=3;
					out<=170;
				end
				if(in == 1) begin
					state<=1;
					out<=171;
				end
				if(in == 2) begin
					state<=10;
					out<=172;
				end
				if(in == 3) begin
					state<=3;
					out<=173;
				end
				if(in == 4) begin
					state<=11;
					out<=174;
				end
				if(in == 5) begin
					state<=3;
					out<=175;
				end
				if(in == 6) begin
					state<=11;
					out<=176;
				end
				if(in == 7) begin
					state<=11;
					out<=177;
				end
				if(in == 8) begin
					state<=11;
					out<=178;
				end
				if(in == 9) begin
					state<=11;
					out<=179;
				end
				if(in == 10) begin
					state<=11;
					out<=180;
				end
				if(in == 11) begin
					state<=11;
					out<=181;
				end
				if(in == 12) begin
					state<=11;
					out<=182;
				end
				if(in == 13) begin
					state<=11;
					out<=183;
				end
				if(in == 14) begin
					state<=11;
					out<=184;
				end
				if(in == 15) begin
					state<=11;
					out<=185;
				end
				if(in == 16) begin
					state<=11;
					out<=186;
				end
				if(in == 17) begin
					state<=11;
					out<=187;
				end
				if(in == 18) begin
					state<=11;
					out<=188;
				end
				if(in == 19) begin
					state<=11;
					out<=189;
				end
				if(in == 20) begin
					state<=11;
					out<=190;
				end
				if(in == 21) begin
					state<=11;
					out<=191;
				end
				if(in == 22) begin
					state<=11;
					out<=192;
				end
				if(in == 23) begin
					state<=11;
					out<=193;
				end
				if(in == 24) begin
					state<=11;
					out<=194;
				end
				if(in == 25) begin
					state<=11;
					out<=195;
				end
				if(in == 26) begin
					state<=11;
					out<=196;
				end
				if(in == 27) begin
					state<=11;
					out<=197;
				end
				if(in == 28) begin
					state<=11;
					out<=198;
				end
				if(in == 29) begin
					state<=11;
					out<=199;
				end
				if(in == 30) begin
					state<=11;
					out<=200;
				end
				if(in == 31) begin
					state<=11;
					out<=201;
				end
				if(in == 32) begin
					state<=11;
					out<=202;
				end
				if(in == 33) begin
					state<=11;
					out<=203;
				end
				if(in == 34) begin
					state<=11;
					out<=204;
				end
				if(in == 35) begin
					state<=11;
					out<=205;
				end
				if(in == 36) begin
					state<=11;
					out<=206;
				end
				if(in == 37) begin
					state<=11;
					out<=207;
				end
				if(in == 38) begin
					state<=11;
					out<=208;
				end
				if(in == 39) begin
					state<=11;
					out<=209;
				end
				if(in == 40) begin
					state<=11;
					out<=210;
				end
				if(in == 41) begin
					state<=11;
					out<=211;
				end
				if(in == 42) begin
					state<=11;
					out<=212;
				end
				if(in == 43) begin
					state<=11;
					out<=213;
				end
				if(in == 44) begin
					state<=11;
					out<=214;
				end
				if(in == 45) begin
					state<=11;
					out<=215;
				end
				if(in == 46) begin
					state<=11;
					out<=216;
				end
				if(in == 47) begin
					state<=11;
					out<=217;
				end
				if(in == 48) begin
					state<=11;
					out<=218;
				end
				if(in == 49) begin
					state<=11;
					out<=219;
				end
				if(in == 50) begin
					state<=11;
					out<=220;
				end
				if(in == 51) begin
					state<=11;
					out<=221;
				end
				if(in == 52) begin
					state<=11;
					out<=222;
				end
				if(in == 53) begin
					state<=3;
					out<=223;
				end
				if(in == 54) begin
					state<=10;
					out<=224;
				end
				if(in == 55) begin
					state<=3;
					out<=225;
				end
				if(in == 56) begin
					state<=11;
					out<=226;
				end
				if(in == 57) begin
					state<=3;
					out<=227;
				end
				if(in == 58) begin
					state<=11;
					out<=228;
				end
				if(in == 59) begin
					state<=11;
					out<=229;
				end
				if(in == 60) begin
					state<=11;
					out<=230;
				end
				if(in == 61) begin
					state<=11;
					out<=231;
				end
				if(in == 62) begin
					state<=11;
					out<=232;
				end
				if(in == 63) begin
					state<=11;
					out<=233;
				end
				if(in == 64) begin
					state<=11;
					out<=234;
				end
				if(in == 65) begin
					state<=11;
					out<=235;
				end
				if(in == 66) begin
					state<=11;
					out<=236;
				end
				if(in == 67) begin
					state<=11;
					out<=237;
				end
				if(in == 68) begin
					state<=11;
					out<=238;
				end
				if(in == 69) begin
					state<=11;
					out<=239;
				end
				if(in == 70) begin
					state<=11;
					out<=240;
				end
				if(in == 71) begin
					state<=11;
					out<=241;
				end
				if(in == 72) begin
					state<=11;
					out<=242;
				end
				if(in == 73) begin
					state<=11;
					out<=243;
				end
				if(in == 74) begin
					state<=11;
					out<=244;
				end
				if(in == 75) begin
					state<=11;
					out<=245;
				end
				if(in == 76) begin
					state<=11;
					out<=246;
				end
				if(in == 77) begin
					state<=11;
					out<=247;
				end
				if(in == 78) begin
					state<=11;
					out<=248;
				end
				if(in == 79) begin
					state<=11;
					out<=249;
				end
				if(in == 80) begin
					state<=11;
					out<=250;
				end
				if(in == 81) begin
					state<=11;
					out<=251;
				end
				if(in == 82) begin
					state<=11;
					out<=252;
				end
				if(in == 83) begin
					state<=11;
					out<=253;
				end
				if(in == 84) begin
					state<=11;
					out<=254;
				end
				if(in == 85) begin
					state<=11;
					out<=255;
				end
				if(in == 86) begin
					state<=11;
					out<=0;
				end
				if(in == 87) begin
					state<=11;
					out<=1;
				end
				if(in == 88) begin
					state<=11;
					out<=2;
				end
				if(in == 89) begin
					state<=11;
					out<=3;
				end
				if(in == 90) begin
					state<=11;
					out<=4;
				end
				if(in == 91) begin
					state<=11;
					out<=5;
				end
				if(in == 92) begin
					state<=11;
					out<=6;
				end
				if(in == 93) begin
					state<=11;
					out<=7;
				end
				if(in == 94) begin
					state<=11;
					out<=8;
				end
				if(in == 95) begin
					state<=11;
					out<=9;
				end
				if(in == 96) begin
					state<=11;
					out<=10;
				end
				if(in == 97) begin
					state<=11;
					out<=11;
				end
				if(in == 98) begin
					state<=11;
					out<=12;
				end
				if(in == 99) begin
					state<=11;
					out<=13;
				end
				if(in == 100) begin
					state<=11;
					out<=14;
				end
				if(in == 101) begin
					state<=11;
					out<=15;
				end
				if(in == 102) begin
					state<=11;
					out<=16;
				end
				if(in == 103) begin
					state<=11;
					out<=17;
				end
				if(in == 104) begin
					state<=11;
					out<=18;
				end
				if(in == 105) begin
					state<=2;
					out<=19;
				end
				if(in == 106) begin
					state<=2;
					out<=20;
				end
				if(in == 107) begin
					state<=2;
					out<=21;
				end
				if(in == 108) begin
					state<=2;
					out<=22;
				end
				if(in == 109) begin
					state<=2;
					out<=23;
				end
				if(in == 110) begin
					state<=2;
					out<=24;
				end
				if(in == 111) begin
					state<=2;
					out<=25;
				end
				if(in == 112) begin
					state<=2;
					out<=26;
				end
				if(in == 113) begin
					state<=2;
					out<=27;
				end
				if(in == 114) begin
					state<=2;
					out<=28;
				end
				if(in == 115) begin
					state<=2;
					out<=29;
				end
				if(in == 116) begin
					state<=2;
					out<=30;
				end
				if(in == 117) begin
					state<=3;
					out<=31;
				end
				if(in == 118) begin
					state<=10;
					out<=32;
				end
				if(in == 119) begin
					state<=3;
					out<=33;
				end
				if(in == 120) begin
					state<=11;
					out<=34;
				end
				if(in == 121) begin
					state<=3;
					out<=35;
				end
				if(in == 122) begin
					state<=11;
					out<=36;
				end
				if(in == 123) begin
					state<=11;
					out<=37;
				end
				if(in == 124) begin
					state<=11;
					out<=38;
				end
				if(in == 125) begin
					state<=11;
					out<=39;
				end
				if(in == 126) begin
					state<=11;
					out<=40;
				end
				if(in == 127) begin
					state<=11;
					out<=41;
				end
				if(in == 128) begin
					state<=11;
					out<=42;
				end
				if(in == 129) begin
					state<=11;
					out<=43;
				end
				if(in == 130) begin
					state<=11;
					out<=44;
				end
				if(in == 131) begin
					state<=11;
					out<=45;
				end
				if(in == 132) begin
					state<=11;
					out<=46;
				end
				if(in == 133) begin
					state<=11;
					out<=47;
				end
				if(in == 134) begin
					state<=11;
					out<=48;
				end
				if(in == 135) begin
					state<=11;
					out<=49;
				end
				if(in == 136) begin
					state<=11;
					out<=50;
				end
				if(in == 137) begin
					state<=11;
					out<=51;
				end
				if(in == 138) begin
					state<=11;
					out<=52;
				end
				if(in == 139) begin
					state<=11;
					out<=53;
				end
				if(in == 140) begin
					state<=11;
					out<=54;
				end
				if(in == 141) begin
					state<=11;
					out<=55;
				end
				if(in == 142) begin
					state<=11;
					out<=56;
				end
				if(in == 143) begin
					state<=11;
					out<=57;
				end
				if(in == 144) begin
					state<=11;
					out<=58;
				end
				if(in == 145) begin
					state<=11;
					out<=59;
				end
				if(in == 146) begin
					state<=11;
					out<=60;
				end
				if(in == 147) begin
					state<=11;
					out<=61;
				end
				if(in == 148) begin
					state<=11;
					out<=62;
				end
				if(in == 149) begin
					state<=11;
					out<=63;
				end
				if(in == 150) begin
					state<=11;
					out<=64;
				end
				if(in == 151) begin
					state<=11;
					out<=65;
				end
				if(in == 152) begin
					state<=11;
					out<=66;
				end
				if(in == 153) begin
					state<=11;
					out<=67;
				end
				if(in == 154) begin
					state<=11;
					out<=68;
				end
				if(in == 155) begin
					state<=11;
					out<=69;
				end
				if(in == 156) begin
					state<=11;
					out<=70;
				end
				if(in == 157) begin
					state<=11;
					out<=71;
				end
				if(in == 158) begin
					state<=11;
					out<=72;
				end
				if(in == 159) begin
					state<=11;
					out<=73;
				end
				if(in == 160) begin
					state<=11;
					out<=74;
				end
				if(in == 161) begin
					state<=11;
					out<=75;
				end
				if(in == 162) begin
					state<=11;
					out<=76;
				end
				if(in == 163) begin
					state<=11;
					out<=77;
				end
				if(in == 164) begin
					state<=11;
					out<=78;
				end
				if(in == 165) begin
					state<=11;
					out<=79;
				end
				if(in == 166) begin
					state<=11;
					out<=80;
				end
				if(in == 167) begin
					state<=11;
					out<=81;
				end
				if(in == 168) begin
					state<=11;
					out<=82;
				end
				if(in == 169) begin
					state<=3;
					out<=83;
				end
				if(in == 170) begin
					state<=10;
					out<=84;
				end
				if(in == 171) begin
					state<=3;
					out<=85;
				end
				if(in == 172) begin
					state<=11;
					out<=86;
				end
				if(in == 173) begin
					state<=3;
					out<=87;
				end
				if(in == 174) begin
					state<=11;
					out<=88;
				end
				if(in == 175) begin
					state<=11;
					out<=89;
				end
				if(in == 176) begin
					state<=11;
					out<=90;
				end
				if(in == 177) begin
					state<=11;
					out<=91;
				end
				if(in == 178) begin
					state<=11;
					out<=92;
				end
				if(in == 179) begin
					state<=11;
					out<=93;
				end
				if(in == 180) begin
					state<=11;
					out<=94;
				end
				if(in == 181) begin
					state<=11;
					out<=95;
				end
				if(in == 182) begin
					state<=11;
					out<=96;
				end
				if(in == 183) begin
					state<=11;
					out<=97;
				end
				if(in == 184) begin
					state<=11;
					out<=98;
				end
				if(in == 185) begin
					state<=11;
					out<=99;
				end
				if(in == 186) begin
					state<=11;
					out<=100;
				end
				if(in == 187) begin
					state<=11;
					out<=101;
				end
				if(in == 188) begin
					state<=11;
					out<=102;
				end
				if(in == 189) begin
					state<=11;
					out<=103;
				end
				if(in == 190) begin
					state<=11;
					out<=104;
				end
				if(in == 191) begin
					state<=11;
					out<=105;
				end
				if(in == 192) begin
					state<=11;
					out<=106;
				end
				if(in == 193) begin
					state<=11;
					out<=107;
				end
				if(in == 194) begin
					state<=11;
					out<=108;
				end
				if(in == 195) begin
					state<=11;
					out<=109;
				end
				if(in == 196) begin
					state<=11;
					out<=110;
				end
				if(in == 197) begin
					state<=11;
					out<=111;
				end
				if(in == 198) begin
					state<=11;
					out<=112;
				end
				if(in == 199) begin
					state<=11;
					out<=113;
				end
				if(in == 200) begin
					state<=11;
					out<=114;
				end
				if(in == 201) begin
					state<=11;
					out<=115;
				end
				if(in == 202) begin
					state<=11;
					out<=116;
				end
				if(in == 203) begin
					state<=11;
					out<=117;
				end
				if(in == 204) begin
					state<=11;
					out<=118;
				end
				if(in == 205) begin
					state<=11;
					out<=119;
				end
				if(in == 206) begin
					state<=11;
					out<=120;
				end
				if(in == 207) begin
					state<=11;
					out<=121;
				end
				if(in == 208) begin
					state<=11;
					out<=122;
				end
				if(in == 209) begin
					state<=11;
					out<=123;
				end
				if(in == 210) begin
					state<=11;
					out<=124;
				end
				if(in == 211) begin
					state<=11;
					out<=125;
				end
				if(in == 212) begin
					state<=11;
					out<=126;
				end
				if(in == 213) begin
					state<=11;
					out<=127;
				end
				if(in == 214) begin
					state<=11;
					out<=128;
				end
				if(in == 215) begin
					state<=11;
					out<=129;
				end
				if(in == 216) begin
					state<=11;
					out<=130;
				end
				if(in == 217) begin
					state<=11;
					out<=131;
				end
				if(in == 218) begin
					state<=11;
					out<=132;
				end
				if(in == 219) begin
					state<=11;
					out<=133;
				end
				if(in == 220) begin
					state<=11;
					out<=134;
				end
				if(in == 221) begin
					state<=2;
					out<=135;
				end
				if(in == 222) begin
					state<=2;
					out<=136;
				end
				if(in == 223) begin
					state<=2;
					out<=137;
				end
				if(in == 224) begin
					state<=2;
					out<=138;
				end
				if(in == 225) begin
					state<=2;
					out<=139;
				end
				if(in == 226) begin
					state<=2;
					out<=140;
				end
				if(in == 227) begin
					state<=2;
					out<=141;
				end
				if(in == 228) begin
					state<=2;
					out<=142;
				end
				if(in == 229) begin
					state<=2;
					out<=143;
				end
				if(in == 230) begin
					state<=2;
					out<=144;
				end
				if(in == 231) begin
					state<=2;
					out<=145;
				end
				if(in == 232) begin
					state<=2;
					out<=146;
				end
				if(in == 233) begin
					state<=3;
					out<=147;
				end
				if(in == 234) begin
					state<=10;
					out<=148;
				end
				if(in == 235) begin
					state<=3;
					out<=149;
				end
				if(in == 236) begin
					state<=11;
					out<=150;
				end
				if(in == 237) begin
					state<=3;
					out<=151;
				end
				if(in == 238) begin
					state<=11;
					out<=152;
				end
				if(in == 239) begin
					state<=11;
					out<=153;
				end
				if(in == 240) begin
					state<=11;
					out<=154;
				end
				if(in == 241) begin
					state<=11;
					out<=155;
				end
				if(in == 242) begin
					state<=11;
					out<=156;
				end
				if(in == 243) begin
					state<=11;
					out<=157;
				end
				if(in == 244) begin
					state<=11;
					out<=158;
				end
				if(in == 245) begin
					state<=11;
					out<=159;
				end
				if(in == 246) begin
					state<=11;
					out<=160;
				end
				if(in == 247) begin
					state<=11;
					out<=161;
				end
				if(in == 248) begin
					state<=11;
					out<=162;
				end
				if(in == 249) begin
					state<=11;
					out<=163;
				end
				if(in == 250) begin
					state<=11;
					out<=164;
				end
				if(in == 251) begin
					state<=11;
					out<=165;
				end
				if(in == 252) begin
					state<=11;
					out<=166;
				end
				if(in == 253) begin
					state<=11;
					out<=167;
				end
				if(in == 254) begin
					state<=11;
					out<=168;
				end
				if(in == 255) begin
					state<=11;
					out<=169;
				end
				if(in == 256) begin
					state<=11;
					out<=170;
				end
				if(in == 257) begin
					state<=11;
					out<=171;
				end
				if(in == 258) begin
					state<=11;
					out<=172;
				end
				if(in == 259) begin
					state<=11;
					out<=173;
				end
				if(in == 260) begin
					state<=11;
					out<=174;
				end
				if(in == 261) begin
					state<=11;
					out<=175;
				end
				if(in == 262) begin
					state<=11;
					out<=176;
				end
				if(in == 263) begin
					state<=11;
					out<=177;
				end
				if(in == 264) begin
					state<=11;
					out<=178;
				end
				if(in == 265) begin
					state<=11;
					out<=179;
				end
				if(in == 266) begin
					state<=11;
					out<=180;
				end
				if(in == 267) begin
					state<=11;
					out<=181;
				end
				if(in == 268) begin
					state<=11;
					out<=182;
				end
				if(in == 269) begin
					state<=11;
					out<=183;
				end
				if(in == 270) begin
					state<=11;
					out<=184;
				end
				if(in == 271) begin
					state<=11;
					out<=185;
				end
				if(in == 272) begin
					state<=11;
					out<=186;
				end
				if(in == 273) begin
					state<=11;
					out<=187;
				end
				if(in == 274) begin
					state<=11;
					out<=188;
				end
				if(in == 275) begin
					state<=11;
					out<=189;
				end
				if(in == 276) begin
					state<=11;
					out<=190;
				end
				if(in == 277) begin
					state<=11;
					out<=191;
				end
				if(in == 278) begin
					state<=11;
					out<=192;
				end
				if(in == 279) begin
					state<=11;
					out<=193;
				end
				if(in == 280) begin
					state<=11;
					out<=194;
				end
				if(in == 281) begin
					state<=11;
					out<=195;
				end
				if(in == 282) begin
					state<=11;
					out<=196;
				end
				if(in == 283) begin
					state<=11;
					out<=197;
				end
				if(in == 284) begin
					state<=11;
					out<=198;
				end
				if(in == 285) begin
					state<=3;
					out<=199;
				end
				if(in == 286) begin
					state<=10;
					out<=200;
				end
				if(in == 287) begin
					state<=3;
					out<=201;
				end
				if(in == 288) begin
					state<=11;
					out<=202;
				end
				if(in == 289) begin
					state<=3;
					out<=203;
				end
				if(in == 290) begin
					state<=11;
					out<=204;
				end
				if(in == 291) begin
					state<=11;
					out<=205;
				end
				if(in == 292) begin
					state<=11;
					out<=206;
				end
				if(in == 293) begin
					state<=11;
					out<=207;
				end
				if(in == 294) begin
					state<=11;
					out<=208;
				end
				if(in == 295) begin
					state<=11;
					out<=209;
				end
				if(in == 296) begin
					state<=11;
					out<=210;
				end
				if(in == 297) begin
					state<=11;
					out<=211;
				end
				if(in == 298) begin
					state<=11;
					out<=212;
				end
				if(in == 299) begin
					state<=11;
					out<=213;
				end
				if(in == 300) begin
					state<=11;
					out<=214;
				end
				if(in == 301) begin
					state<=11;
					out<=215;
				end
				if(in == 302) begin
					state<=11;
					out<=216;
				end
				if(in == 303) begin
					state<=11;
					out<=217;
				end
				if(in == 304) begin
					state<=11;
					out<=218;
				end
				if(in == 305) begin
					state<=11;
					out<=219;
				end
				if(in == 306) begin
					state<=11;
					out<=220;
				end
				if(in == 307) begin
					state<=11;
					out<=221;
				end
				if(in == 308) begin
					state<=11;
					out<=222;
				end
				if(in == 309) begin
					state<=11;
					out<=223;
				end
				if(in == 310) begin
					state<=11;
					out<=224;
				end
				if(in == 311) begin
					state<=11;
					out<=225;
				end
				if(in == 312) begin
					state<=11;
					out<=226;
				end
				if(in == 313) begin
					state<=11;
					out<=227;
				end
				if(in == 314) begin
					state<=11;
					out<=228;
				end
				if(in == 315) begin
					state<=11;
					out<=229;
				end
				if(in == 316) begin
					state<=11;
					out<=230;
				end
				if(in == 317) begin
					state<=11;
					out<=231;
				end
				if(in == 318) begin
					state<=11;
					out<=232;
				end
				if(in == 319) begin
					state<=11;
					out<=233;
				end
				if(in == 320) begin
					state<=11;
					out<=234;
				end
				if(in == 321) begin
					state<=11;
					out<=235;
				end
				if(in == 322) begin
					state<=11;
					out<=236;
				end
				if(in == 323) begin
					state<=11;
					out<=237;
				end
				if(in == 324) begin
					state<=11;
					out<=238;
				end
				if(in == 325) begin
					state<=11;
					out<=239;
				end
				if(in == 326) begin
					state<=11;
					out<=240;
				end
				if(in == 327) begin
					state<=11;
					out<=241;
				end
				if(in == 328) begin
					state<=11;
					out<=242;
				end
				if(in == 329) begin
					state<=11;
					out<=243;
				end
				if(in == 330) begin
					state<=11;
					out<=244;
				end
				if(in == 331) begin
					state<=11;
					out<=245;
				end
				if(in == 332) begin
					state<=11;
					out<=246;
				end
				if(in == 333) begin
					state<=11;
					out<=247;
				end
				if(in == 334) begin
					state<=11;
					out<=248;
				end
				if(in == 335) begin
					state<=11;
					out<=249;
				end
				if(in == 336) begin
					state<=11;
					out<=250;
				end
				if(in == 337) begin
					state<=2;
					out<=251;
				end
				if(in == 338) begin
					state<=2;
					out<=252;
				end
				if(in == 339) begin
					state<=2;
					out<=253;
				end
				if(in == 340) begin
					state<=2;
					out<=254;
				end
				if(in == 341) begin
					state<=2;
					out<=255;
				end
				if(in == 342) begin
					state<=2;
					out<=0;
				end
				if(in == 343) begin
					state<=2;
					out<=1;
				end
				if(in == 344) begin
					state<=2;
					out<=2;
				end
				if(in == 345) begin
					state<=2;
					out<=3;
				end
				if(in == 346) begin
					state<=2;
					out<=4;
				end
				if(in == 347) begin
					state<=2;
					out<=5;
				end
				if(in == 348) begin
					state<=2;
					out<=6;
				end
				if(in == 349) begin
					state<=3;
					out<=7;
				end
				if(in == 350) begin
					state<=10;
					out<=8;
				end
				if(in == 351) begin
					state<=3;
					out<=9;
				end
				if(in == 352) begin
					state<=11;
					out<=10;
				end
				if(in == 353) begin
					state<=3;
					out<=11;
				end
				if(in == 354) begin
					state<=11;
					out<=12;
				end
				if(in == 355) begin
					state<=11;
					out<=13;
				end
				if(in == 356) begin
					state<=11;
					out<=14;
				end
				if(in == 357) begin
					state<=11;
					out<=15;
				end
				if(in == 358) begin
					state<=11;
					out<=16;
				end
				if(in == 359) begin
					state<=11;
					out<=17;
				end
				if(in == 360) begin
					state<=11;
					out<=18;
				end
				if(in == 361) begin
					state<=11;
					out<=19;
				end
				if(in == 362) begin
					state<=11;
					out<=20;
				end
				if(in == 363) begin
					state<=11;
					out<=21;
				end
				if(in == 364) begin
					state<=11;
					out<=22;
				end
				if(in == 365) begin
					state<=11;
					out<=23;
				end
				if(in == 366) begin
					state<=11;
					out<=24;
				end
				if(in == 367) begin
					state<=11;
					out<=25;
				end
				if(in == 368) begin
					state<=11;
					out<=26;
				end
				if(in == 369) begin
					state<=11;
					out<=27;
				end
				if(in == 370) begin
					state<=11;
					out<=28;
				end
				if(in == 371) begin
					state<=11;
					out<=29;
				end
				if(in == 372) begin
					state<=11;
					out<=30;
				end
				if(in == 373) begin
					state<=11;
					out<=31;
				end
				if(in == 374) begin
					state<=11;
					out<=32;
				end
				if(in == 375) begin
					state<=11;
					out<=33;
				end
				if(in == 376) begin
					state<=11;
					out<=34;
				end
				if(in == 377) begin
					state<=11;
					out<=35;
				end
				if(in == 378) begin
					state<=11;
					out<=36;
				end
				if(in == 379) begin
					state<=11;
					out<=37;
				end
				if(in == 380) begin
					state<=11;
					out<=38;
				end
				if(in == 381) begin
					state<=11;
					out<=39;
				end
				if(in == 382) begin
					state<=11;
					out<=40;
				end
				if(in == 383) begin
					state<=11;
					out<=41;
				end
				if(in == 384) begin
					state<=11;
					out<=42;
				end
				if(in == 385) begin
					state<=11;
					out<=43;
				end
				if(in == 386) begin
					state<=11;
					out<=44;
				end
				if(in == 387) begin
					state<=11;
					out<=45;
				end
				if(in == 388) begin
					state<=11;
					out<=46;
				end
				if(in == 389) begin
					state<=11;
					out<=47;
				end
				if(in == 390) begin
					state<=11;
					out<=48;
				end
				if(in == 391) begin
					state<=11;
					out<=49;
				end
				if(in == 392) begin
					state<=11;
					out<=50;
				end
				if(in == 393) begin
					state<=11;
					out<=51;
				end
				if(in == 394) begin
					state<=11;
					out<=52;
				end
				if(in == 395) begin
					state<=11;
					out<=53;
				end
				if(in == 396) begin
					state<=11;
					out<=54;
				end
				if(in == 397) begin
					state<=11;
					out<=55;
				end
				if(in == 398) begin
					state<=11;
					out<=56;
				end
				if(in == 399) begin
					state<=11;
					out<=57;
				end
				if(in == 400) begin
					state<=11;
					out<=58;
				end
				if(in == 401) begin
					state<=3;
					out<=59;
				end
				if(in == 402) begin
					state<=10;
					out<=60;
				end
				if(in == 403) begin
					state<=3;
					out<=61;
				end
				if(in == 404) begin
					state<=11;
					out<=62;
				end
				if(in == 405) begin
					state<=3;
					out<=63;
				end
				if(in == 406) begin
					state<=11;
					out<=64;
				end
				if(in == 407) begin
					state<=11;
					out<=65;
				end
				if(in == 408) begin
					state<=11;
					out<=66;
				end
				if(in == 409) begin
					state<=11;
					out<=67;
				end
				if(in == 410) begin
					state<=11;
					out<=68;
				end
				if(in == 411) begin
					state<=11;
					out<=69;
				end
				if(in == 412) begin
					state<=11;
					out<=70;
				end
				if(in == 413) begin
					state<=11;
					out<=71;
				end
				if(in == 414) begin
					state<=11;
					out<=72;
				end
				if(in == 415) begin
					state<=11;
					out<=73;
				end
				if(in == 416) begin
					state<=11;
					out<=74;
				end
				if(in == 417) begin
					state<=11;
					out<=75;
				end
				if(in == 418) begin
					state<=11;
					out<=76;
				end
				if(in == 419) begin
					state<=11;
					out<=77;
				end
				if(in == 420) begin
					state<=11;
					out<=78;
				end
				if(in == 421) begin
					state<=11;
					out<=79;
				end
				if(in == 422) begin
					state<=11;
					out<=80;
				end
				if(in == 423) begin
					state<=11;
					out<=81;
				end
				if(in == 424) begin
					state<=11;
					out<=82;
				end
				if(in == 425) begin
					state<=11;
					out<=83;
				end
				if(in == 426) begin
					state<=11;
					out<=84;
				end
				if(in == 427) begin
					state<=11;
					out<=85;
				end
				if(in == 428) begin
					state<=11;
					out<=86;
				end
				if(in == 429) begin
					state<=11;
					out<=87;
				end
				if(in == 430) begin
					state<=11;
					out<=88;
				end
				if(in == 431) begin
					state<=11;
					out<=89;
				end
				if(in == 432) begin
					state<=11;
					out<=90;
				end
				if(in == 433) begin
					state<=11;
					out<=91;
				end
				if(in == 434) begin
					state<=11;
					out<=92;
				end
				if(in == 435) begin
					state<=11;
					out<=93;
				end
				if(in == 436) begin
					state<=11;
					out<=94;
				end
				if(in == 437) begin
					state<=11;
					out<=95;
				end
				if(in == 438) begin
					state<=11;
					out<=96;
				end
				if(in == 439) begin
					state<=11;
					out<=97;
				end
				if(in == 440) begin
					state<=11;
					out<=98;
				end
				if(in == 441) begin
					state<=11;
					out<=99;
				end
				if(in == 442) begin
					state<=11;
					out<=100;
				end
				if(in == 443) begin
					state<=11;
					out<=101;
				end
				if(in == 444) begin
					state<=11;
					out<=102;
				end
				if(in == 445) begin
					state<=11;
					out<=103;
				end
				if(in == 446) begin
					state<=11;
					out<=104;
				end
				if(in == 447) begin
					state<=11;
					out<=105;
				end
				if(in == 448) begin
					state<=11;
					out<=106;
				end
				if(in == 449) begin
					state<=11;
					out<=107;
				end
				if(in == 450) begin
					state<=11;
					out<=108;
				end
				if(in == 451) begin
					state<=11;
					out<=109;
				end
				if(in == 452) begin
					state<=11;
					out<=110;
				end
				if(in == 453) begin
					state<=2;
					out<=111;
				end
				if(in == 454) begin
					state<=2;
					out<=112;
				end
				if(in == 455) begin
					state<=2;
					out<=113;
				end
				if(in == 456) begin
					state<=2;
					out<=114;
				end
				if(in == 457) begin
					state<=2;
					out<=115;
				end
				if(in == 458) begin
					state<=2;
					out<=116;
				end
				if(in == 459) begin
					state<=2;
					out<=117;
				end
				if(in == 460) begin
					state<=2;
					out<=118;
				end
				if(in == 461) begin
					state<=2;
					out<=119;
				end
				if(in == 462) begin
					state<=2;
					out<=120;
				end
				if(in == 463) begin
					state<=2;
					out<=121;
				end
				if(in == 464) begin
					state<=2;
					out<=122;
				end
				if(in == 465) begin
					state<=3;
					out<=123;
				end
				if(in == 466) begin
					state<=10;
					out<=124;
				end
				if(in == 467) begin
					state<=3;
					out<=125;
				end
				if(in == 468) begin
					state<=11;
					out<=126;
				end
				if(in == 469) begin
					state<=3;
					out<=127;
				end
				if(in == 470) begin
					state<=11;
					out<=128;
				end
				if(in == 471) begin
					state<=11;
					out<=129;
				end
				if(in == 472) begin
					state<=11;
					out<=130;
				end
				if(in == 473) begin
					state<=11;
					out<=131;
				end
				if(in == 474) begin
					state<=11;
					out<=132;
				end
				if(in == 475) begin
					state<=11;
					out<=133;
				end
				if(in == 476) begin
					state<=11;
					out<=134;
				end
				if(in == 477) begin
					state<=11;
					out<=135;
				end
				if(in == 478) begin
					state<=11;
					out<=136;
				end
				if(in == 479) begin
					state<=11;
					out<=137;
				end
				if(in == 480) begin
					state<=11;
					out<=138;
				end
				if(in == 481) begin
					state<=11;
					out<=139;
				end
				if(in == 482) begin
					state<=11;
					out<=140;
				end
				if(in == 483) begin
					state<=11;
					out<=141;
				end
				if(in == 484) begin
					state<=11;
					out<=142;
				end
				if(in == 485) begin
					state<=11;
					out<=143;
				end
				if(in == 486) begin
					state<=11;
					out<=144;
				end
				if(in == 487) begin
					state<=11;
					out<=145;
				end
				if(in == 488) begin
					state<=11;
					out<=146;
				end
				if(in == 489) begin
					state<=11;
					out<=147;
				end
				if(in == 490) begin
					state<=11;
					out<=148;
				end
				if(in == 491) begin
					state<=11;
					out<=149;
				end
				if(in == 492) begin
					state<=11;
					out<=150;
				end
				if(in == 493) begin
					state<=11;
					out<=151;
				end
				if(in == 494) begin
					state<=11;
					out<=152;
				end
				if(in == 495) begin
					state<=11;
					out<=153;
				end
				if(in == 496) begin
					state<=11;
					out<=154;
				end
				if(in == 497) begin
					state<=11;
					out<=155;
				end
				if(in == 498) begin
					state<=11;
					out<=156;
				end
				if(in == 499) begin
					state<=11;
					out<=157;
				end
				if(in == 500) begin
					state<=11;
					out<=158;
				end
				if(in == 501) begin
					state<=11;
					out<=159;
				end
				if(in == 502) begin
					state<=11;
					out<=160;
				end
				if(in == 503) begin
					state<=11;
					out<=161;
				end
				if(in == 504) begin
					state<=11;
					out<=162;
				end
				if(in == 505) begin
					state<=11;
					out<=163;
				end
				if(in == 506) begin
					state<=11;
					out<=164;
				end
				if(in == 507) begin
					state<=11;
					out<=165;
				end
				if(in == 508) begin
					state<=11;
					out<=166;
				end
				if(in == 509) begin
					state<=11;
					out<=167;
				end
				if(in == 510) begin
					state<=11;
					out<=168;
				end
				if(in == 511) begin
					state<=11;
					out<=169;
				end
				if(in == 512) begin
					state<=11;
					out<=170;
				end
				if(in == 513) begin
					state<=11;
					out<=171;
				end
				if(in == 514) begin
					state<=11;
					out<=172;
				end
				if(in == 515) begin
					state<=11;
					out<=173;
				end
				if(in == 516) begin
					state<=11;
					out<=174;
				end
				if(in == 517) begin
					state<=3;
					out<=175;
				end
				if(in == 518) begin
					state<=10;
					out<=176;
				end
				if(in == 519) begin
					state<=3;
					out<=177;
				end
				if(in == 520) begin
					state<=11;
					out<=178;
				end
				if(in == 521) begin
					state<=3;
					out<=179;
				end
				if(in == 522) begin
					state<=11;
					out<=180;
				end
				if(in == 523) begin
					state<=11;
					out<=181;
				end
				if(in == 524) begin
					state<=11;
					out<=182;
				end
				if(in == 525) begin
					state<=11;
					out<=183;
				end
				if(in == 526) begin
					state<=11;
					out<=184;
				end
				if(in == 527) begin
					state<=11;
					out<=185;
				end
				if(in == 528) begin
					state<=11;
					out<=186;
				end
				if(in == 529) begin
					state<=11;
					out<=187;
				end
				if(in == 530) begin
					state<=11;
					out<=188;
				end
				if(in == 531) begin
					state<=11;
					out<=189;
				end
				if(in == 532) begin
					state<=11;
					out<=190;
				end
				if(in == 533) begin
					state<=11;
					out<=191;
				end
				if(in == 534) begin
					state<=11;
					out<=192;
				end
				if(in == 535) begin
					state<=11;
					out<=193;
				end
				if(in == 536) begin
					state<=11;
					out<=194;
				end
				if(in == 537) begin
					state<=11;
					out<=195;
				end
				if(in == 538) begin
					state<=11;
					out<=196;
				end
				if(in == 539) begin
					state<=11;
					out<=197;
				end
				if(in == 540) begin
					state<=11;
					out<=198;
				end
				if(in == 541) begin
					state<=11;
					out<=199;
				end
				if(in == 542) begin
					state<=11;
					out<=200;
				end
				if(in == 543) begin
					state<=11;
					out<=201;
				end
				if(in == 544) begin
					state<=11;
					out<=202;
				end
				if(in == 545) begin
					state<=11;
					out<=203;
				end
				if(in == 546) begin
					state<=11;
					out<=204;
				end
				if(in == 547) begin
					state<=11;
					out<=205;
				end
				if(in == 548) begin
					state<=11;
					out<=206;
				end
				if(in == 549) begin
					state<=11;
					out<=207;
				end
				if(in == 550) begin
					state<=11;
					out<=208;
				end
				if(in == 551) begin
					state<=11;
					out<=209;
				end
				if(in == 552) begin
					state<=11;
					out<=210;
				end
				if(in == 553) begin
					state<=11;
					out<=211;
				end
				if(in == 554) begin
					state<=11;
					out<=212;
				end
				if(in == 555) begin
					state<=11;
					out<=213;
				end
				if(in == 556) begin
					state<=11;
					out<=214;
				end
				if(in == 557) begin
					state<=11;
					out<=215;
				end
				if(in == 558) begin
					state<=11;
					out<=216;
				end
				if(in == 559) begin
					state<=11;
					out<=217;
				end
				if(in == 560) begin
					state<=11;
					out<=218;
				end
				if(in == 561) begin
					state<=11;
					out<=219;
				end
				if(in == 562) begin
					state<=11;
					out<=220;
				end
				if(in == 563) begin
					state<=11;
					out<=221;
				end
				if(in == 564) begin
					state<=11;
					out<=222;
				end
				if(in == 565) begin
					state<=11;
					out<=223;
				end
				if(in == 566) begin
					state<=11;
					out<=224;
				end
				if(in == 567) begin
					state<=11;
					out<=225;
				end
				if(in == 568) begin
					state<=11;
					out<=226;
				end
				if(in == 569) begin
					state<=2;
					out<=227;
				end
				if(in == 570) begin
					state<=2;
					out<=228;
				end
				if(in == 571) begin
					state<=2;
					out<=229;
				end
				if(in == 572) begin
					state<=2;
					out<=230;
				end
				if(in == 573) begin
					state<=2;
					out<=231;
				end
				if(in == 574) begin
					state<=2;
					out<=232;
				end
				if(in == 575) begin
					state<=2;
					out<=233;
				end
				if(in == 576) begin
					state<=2;
					out<=234;
				end
				if(in == 577) begin
					state<=2;
					out<=235;
				end
				if(in == 578) begin
					state<=2;
					out<=236;
				end
				if(in == 579) begin
					state<=2;
					out<=237;
				end
				if(in == 580) begin
					state<=2;
					out<=238;
				end
				if(in == 581) begin
					state<=3;
					out<=239;
				end
				if(in == 582) begin
					state<=10;
					out<=240;
				end
				if(in == 583) begin
					state<=3;
					out<=241;
				end
				if(in == 584) begin
					state<=11;
					out<=242;
				end
				if(in == 585) begin
					state<=3;
					out<=243;
				end
				if(in == 586) begin
					state<=11;
					out<=244;
				end
				if(in == 587) begin
					state<=11;
					out<=245;
				end
				if(in == 588) begin
					state<=11;
					out<=246;
				end
				if(in == 589) begin
					state<=11;
					out<=247;
				end
				if(in == 590) begin
					state<=11;
					out<=248;
				end
				if(in == 591) begin
					state<=11;
					out<=249;
				end
				if(in == 592) begin
					state<=11;
					out<=250;
				end
				if(in == 593) begin
					state<=11;
					out<=251;
				end
				if(in == 594) begin
					state<=11;
					out<=252;
				end
				if(in == 595) begin
					state<=11;
					out<=253;
				end
				if(in == 596) begin
					state<=11;
					out<=254;
				end
				if(in == 597) begin
					state<=11;
					out<=255;
				end
				if(in == 598) begin
					state<=11;
					out<=0;
				end
				if(in == 599) begin
					state<=11;
					out<=1;
				end
				if(in == 600) begin
					state<=11;
					out<=2;
				end
				if(in == 601) begin
					state<=11;
					out<=3;
				end
				if(in == 602) begin
					state<=11;
					out<=4;
				end
				if(in == 603) begin
					state<=11;
					out<=5;
				end
				if(in == 604) begin
					state<=11;
					out<=6;
				end
				if(in == 605) begin
					state<=11;
					out<=7;
				end
				if(in == 606) begin
					state<=11;
					out<=8;
				end
				if(in == 607) begin
					state<=11;
					out<=9;
				end
				if(in == 608) begin
					state<=11;
					out<=10;
				end
				if(in == 609) begin
					state<=11;
					out<=11;
				end
				if(in == 610) begin
					state<=11;
					out<=12;
				end
				if(in == 611) begin
					state<=11;
					out<=13;
				end
				if(in == 612) begin
					state<=11;
					out<=14;
				end
				if(in == 613) begin
					state<=11;
					out<=15;
				end
				if(in == 614) begin
					state<=11;
					out<=16;
				end
				if(in == 615) begin
					state<=11;
					out<=17;
				end
				if(in == 616) begin
					state<=11;
					out<=18;
				end
				if(in == 617) begin
					state<=11;
					out<=19;
				end
				if(in == 618) begin
					state<=11;
					out<=20;
				end
				if(in == 619) begin
					state<=11;
					out<=21;
				end
				if(in == 620) begin
					state<=11;
					out<=22;
				end
				if(in == 621) begin
					state<=11;
					out<=23;
				end
				if(in == 622) begin
					state<=11;
					out<=24;
				end
				if(in == 623) begin
					state<=11;
					out<=25;
				end
				if(in == 624) begin
					state<=11;
					out<=26;
				end
				if(in == 625) begin
					state<=11;
					out<=27;
				end
				if(in == 626) begin
					state<=11;
					out<=28;
				end
				if(in == 627) begin
					state<=11;
					out<=29;
				end
				if(in == 628) begin
					state<=11;
					out<=30;
				end
				if(in == 629) begin
					state<=11;
					out<=31;
				end
				if(in == 630) begin
					state<=11;
					out<=32;
				end
				if(in == 631) begin
					state<=11;
					out<=33;
				end
				if(in == 632) begin
					state<=11;
					out<=34;
				end
				if(in == 633) begin
					state<=3;
					out<=35;
				end
				if(in == 634) begin
					state<=10;
					out<=36;
				end
				if(in == 635) begin
					state<=3;
					out<=37;
				end
				if(in == 636) begin
					state<=11;
					out<=38;
				end
				if(in == 637) begin
					state<=3;
					out<=39;
				end
				if(in == 638) begin
					state<=11;
					out<=40;
				end
				if(in == 639) begin
					state<=11;
					out<=41;
				end
				if(in == 640) begin
					state<=11;
					out<=42;
				end
				if(in == 641) begin
					state<=11;
					out<=43;
				end
				if(in == 642) begin
					state<=11;
					out<=44;
				end
				if(in == 643) begin
					state<=11;
					out<=45;
				end
				if(in == 644) begin
					state<=11;
					out<=46;
				end
				if(in == 645) begin
					state<=11;
					out<=47;
				end
				if(in == 646) begin
					state<=11;
					out<=48;
				end
				if(in == 647) begin
					state<=11;
					out<=49;
				end
				if(in == 648) begin
					state<=11;
					out<=50;
				end
				if(in == 649) begin
					state<=11;
					out<=51;
				end
				if(in == 650) begin
					state<=11;
					out<=52;
				end
				if(in == 651) begin
					state<=11;
					out<=53;
				end
				if(in == 652) begin
					state<=11;
					out<=54;
				end
				if(in == 653) begin
					state<=11;
					out<=55;
				end
				if(in == 654) begin
					state<=11;
					out<=56;
				end
				if(in == 655) begin
					state<=11;
					out<=57;
				end
				if(in == 656) begin
					state<=11;
					out<=58;
				end
				if(in == 657) begin
					state<=11;
					out<=59;
				end
				if(in == 658) begin
					state<=11;
					out<=60;
				end
				if(in == 659) begin
					state<=11;
					out<=61;
				end
				if(in == 660) begin
					state<=11;
					out<=62;
				end
				if(in == 661) begin
					state<=11;
					out<=63;
				end
				if(in == 662) begin
					state<=11;
					out<=64;
				end
				if(in == 663) begin
					state<=11;
					out<=65;
				end
				if(in == 664) begin
					state<=11;
					out<=66;
				end
				if(in == 665) begin
					state<=11;
					out<=67;
				end
				if(in == 666) begin
					state<=11;
					out<=68;
				end
				if(in == 667) begin
					state<=11;
					out<=69;
				end
				if(in == 668) begin
					state<=11;
					out<=70;
				end
				if(in == 669) begin
					state<=11;
					out<=71;
				end
				if(in == 670) begin
					state<=11;
					out<=72;
				end
				if(in == 671) begin
					state<=11;
					out<=73;
				end
				if(in == 672) begin
					state<=11;
					out<=74;
				end
				if(in == 673) begin
					state<=11;
					out<=75;
				end
				if(in == 674) begin
					state<=11;
					out<=76;
				end
				if(in == 675) begin
					state<=11;
					out<=77;
				end
				if(in == 676) begin
					state<=11;
					out<=78;
				end
				if(in == 677) begin
					state<=11;
					out<=79;
				end
				if(in == 678) begin
					state<=11;
					out<=80;
				end
				if(in == 679) begin
					state<=11;
					out<=81;
				end
				if(in == 680) begin
					state<=11;
					out<=82;
				end
				if(in == 681) begin
					state<=11;
					out<=83;
				end
				if(in == 682) begin
					state<=11;
					out<=84;
				end
				if(in == 683) begin
					state<=11;
					out<=85;
				end
				if(in == 684) begin
					state<=11;
					out<=86;
				end
				if(in == 685) begin
					state<=2;
					out<=87;
				end
				if(in == 686) begin
					state<=2;
					out<=88;
				end
				if(in == 687) begin
					state<=2;
					out<=89;
				end
				if(in == 688) begin
					state<=2;
					out<=90;
				end
				if(in == 689) begin
					state<=2;
					out<=91;
				end
				if(in == 690) begin
					state<=2;
					out<=92;
				end
				if(in == 691) begin
					state<=2;
					out<=93;
				end
				if(in == 692) begin
					state<=2;
					out<=94;
				end
				if(in == 693) begin
					state<=2;
					out<=95;
				end
				if(in == 694) begin
					state<=2;
					out<=96;
				end
				if(in == 695) begin
					state<=2;
					out<=97;
				end
				if(in == 696) begin
					state<=2;
					out<=98;
				end
				if(in == 697) begin
					state<=3;
					out<=99;
				end
				if(in == 698) begin
					state<=10;
					out<=100;
				end
				if(in == 699) begin
					state<=3;
					out<=101;
				end
				if(in == 700) begin
					state<=11;
					out<=102;
				end
				if(in == 701) begin
					state<=3;
					out<=103;
				end
				if(in == 702) begin
					state<=11;
					out<=104;
				end
				if(in == 703) begin
					state<=11;
					out<=105;
				end
				if(in == 704) begin
					state<=11;
					out<=106;
				end
				if(in == 705) begin
					state<=11;
					out<=107;
				end
				if(in == 706) begin
					state<=11;
					out<=108;
				end
				if(in == 707) begin
					state<=11;
					out<=109;
				end
				if(in == 708) begin
					state<=11;
					out<=110;
				end
				if(in == 709) begin
					state<=11;
					out<=111;
				end
				if(in == 710) begin
					state<=11;
					out<=112;
				end
				if(in == 711) begin
					state<=11;
					out<=113;
				end
				if(in == 712) begin
					state<=11;
					out<=114;
				end
				if(in == 713) begin
					state<=11;
					out<=115;
				end
				if(in == 714) begin
					state<=11;
					out<=116;
				end
				if(in == 715) begin
					state<=11;
					out<=117;
				end
				if(in == 716) begin
					state<=11;
					out<=118;
				end
				if(in == 717) begin
					state<=11;
					out<=119;
				end
				if(in == 718) begin
					state<=11;
					out<=120;
				end
				if(in == 719) begin
					state<=11;
					out<=121;
				end
				if(in == 720) begin
					state<=11;
					out<=122;
				end
				if(in == 721) begin
					state<=11;
					out<=123;
				end
				if(in == 722) begin
					state<=11;
					out<=124;
				end
				if(in == 723) begin
					state<=11;
					out<=125;
				end
				if(in == 724) begin
					state<=11;
					out<=126;
				end
				if(in == 725) begin
					state<=11;
					out<=127;
				end
				if(in == 726) begin
					state<=11;
					out<=128;
				end
				if(in == 727) begin
					state<=11;
					out<=129;
				end
				if(in == 728) begin
					state<=11;
					out<=130;
				end
				if(in == 729) begin
					state<=11;
					out<=131;
				end
				if(in == 730) begin
					state<=11;
					out<=132;
				end
				if(in == 731) begin
					state<=11;
					out<=133;
				end
				if(in == 732) begin
					state<=11;
					out<=134;
				end
				if(in == 733) begin
					state<=11;
					out<=135;
				end
				if(in == 734) begin
					state<=11;
					out<=136;
				end
				if(in == 735) begin
					state<=11;
					out<=137;
				end
				if(in == 736) begin
					state<=11;
					out<=138;
				end
				if(in == 737) begin
					state<=11;
					out<=139;
				end
				if(in == 738) begin
					state<=11;
					out<=140;
				end
				if(in == 739) begin
					state<=11;
					out<=141;
				end
				if(in == 740) begin
					state<=11;
					out<=142;
				end
				if(in == 741) begin
					state<=11;
					out<=143;
				end
				if(in == 742) begin
					state<=11;
					out<=144;
				end
				if(in == 743) begin
					state<=11;
					out<=145;
				end
				if(in == 744) begin
					state<=11;
					out<=146;
				end
				if(in == 745) begin
					state<=11;
					out<=147;
				end
				if(in == 746) begin
					state<=11;
					out<=148;
				end
				if(in == 747) begin
					state<=11;
					out<=149;
				end
				if(in == 748) begin
					state<=11;
					out<=150;
				end
				if(in == 749) begin
					state<=3;
					out<=151;
				end
				if(in == 750) begin
					state<=10;
					out<=152;
				end
				if(in == 751) begin
					state<=3;
					out<=153;
				end
				if(in == 752) begin
					state<=11;
					out<=154;
				end
				if(in == 753) begin
					state<=3;
					out<=155;
				end
				if(in == 754) begin
					state<=11;
					out<=156;
				end
				if(in == 755) begin
					state<=11;
					out<=157;
				end
				if(in == 756) begin
					state<=11;
					out<=158;
				end
				if(in == 757) begin
					state<=11;
					out<=159;
				end
				if(in == 758) begin
					state<=11;
					out<=160;
				end
				if(in == 759) begin
					state<=11;
					out<=161;
				end
				if(in == 760) begin
					state<=11;
					out<=162;
				end
				if(in == 761) begin
					state<=11;
					out<=163;
				end
				if(in == 762) begin
					state<=11;
					out<=164;
				end
				if(in == 763) begin
					state<=11;
					out<=165;
				end
				if(in == 764) begin
					state<=11;
					out<=166;
				end
				if(in == 765) begin
					state<=11;
					out<=167;
				end
				if(in == 766) begin
					state<=11;
					out<=168;
				end
				if(in == 767) begin
					state<=11;
					out<=169;
				end
				if(in == 768) begin
					state<=11;
					out<=170;
				end
				if(in == 769) begin
					state<=11;
					out<=171;
				end
				if(in == 770) begin
					state<=11;
					out<=172;
				end
				if(in == 771) begin
					state<=11;
					out<=173;
				end
				if(in == 772) begin
					state<=11;
					out<=174;
				end
				if(in == 773) begin
					state<=11;
					out<=175;
				end
				if(in == 774) begin
					state<=11;
					out<=176;
				end
				if(in == 775) begin
					state<=11;
					out<=177;
				end
				if(in == 776) begin
					state<=11;
					out<=178;
				end
				if(in == 777) begin
					state<=11;
					out<=179;
				end
				if(in == 778) begin
					state<=11;
					out<=180;
				end
				if(in == 779) begin
					state<=11;
					out<=181;
				end
				if(in == 780) begin
					state<=11;
					out<=182;
				end
				if(in == 781) begin
					state<=11;
					out<=183;
				end
				if(in == 782) begin
					state<=11;
					out<=184;
				end
				if(in == 783) begin
					state<=11;
					out<=185;
				end
				if(in == 784) begin
					state<=11;
					out<=186;
				end
				if(in == 785) begin
					state<=11;
					out<=187;
				end
				if(in == 786) begin
					state<=11;
					out<=188;
				end
				if(in == 787) begin
					state<=11;
					out<=189;
				end
				if(in == 788) begin
					state<=11;
					out<=190;
				end
				if(in == 789) begin
					state<=11;
					out<=191;
				end
				if(in == 790) begin
					state<=11;
					out<=192;
				end
				if(in == 791) begin
					state<=11;
					out<=193;
				end
				if(in == 792) begin
					state<=11;
					out<=194;
				end
				if(in == 793) begin
					state<=11;
					out<=195;
				end
				if(in == 794) begin
					state<=11;
					out<=196;
				end
				if(in == 795) begin
					state<=11;
					out<=197;
				end
				if(in == 796) begin
					state<=11;
					out<=198;
				end
				if(in == 797) begin
					state<=11;
					out<=199;
				end
				if(in == 798) begin
					state<=11;
					out<=200;
				end
				if(in == 799) begin
					state<=11;
					out<=201;
				end
				if(in == 800) begin
					state<=11;
					out<=202;
				end
				if(in == 801) begin
					state<=2;
					out<=203;
				end
				if(in == 802) begin
					state<=2;
					out<=204;
				end
				if(in == 803) begin
					state<=2;
					out<=205;
				end
				if(in == 804) begin
					state<=2;
					out<=206;
				end
				if(in == 805) begin
					state<=2;
					out<=207;
				end
				if(in == 806) begin
					state<=2;
					out<=208;
				end
				if(in == 807) begin
					state<=2;
					out<=209;
				end
				if(in == 808) begin
					state<=2;
					out<=210;
				end
				if(in == 809) begin
					state<=2;
					out<=211;
				end
				if(in == 810) begin
					state<=2;
					out<=212;
				end
				if(in == 811) begin
					state<=2;
					out<=213;
				end
				if(in == 812) begin
					state<=2;
					out<=214;
				end
				if(in == 813) begin
					state<=3;
					out<=215;
				end
				if(in == 814) begin
					state<=10;
					out<=216;
				end
				if(in == 815) begin
					state<=3;
					out<=217;
				end
				if(in == 816) begin
					state<=11;
					out<=218;
				end
				if(in == 817) begin
					state<=3;
					out<=219;
				end
				if(in == 818) begin
					state<=11;
					out<=220;
				end
				if(in == 819) begin
					state<=11;
					out<=221;
				end
				if(in == 820) begin
					state<=11;
					out<=222;
				end
				if(in == 821) begin
					state<=11;
					out<=223;
				end
				if(in == 822) begin
					state<=11;
					out<=224;
				end
				if(in == 823) begin
					state<=11;
					out<=225;
				end
				if(in == 824) begin
					state<=11;
					out<=226;
				end
				if(in == 825) begin
					state<=11;
					out<=227;
				end
				if(in == 826) begin
					state<=11;
					out<=228;
				end
				if(in == 827) begin
					state<=11;
					out<=229;
				end
				if(in == 828) begin
					state<=11;
					out<=230;
				end
				if(in == 829) begin
					state<=11;
					out<=231;
				end
				if(in == 830) begin
					state<=11;
					out<=232;
				end
				if(in == 831) begin
					state<=11;
					out<=233;
				end
				if(in == 832) begin
					state<=11;
					out<=234;
				end
				if(in == 833) begin
					state<=11;
					out<=235;
				end
				if(in == 834) begin
					state<=11;
					out<=236;
				end
				if(in == 835) begin
					state<=11;
					out<=237;
				end
				if(in == 836) begin
					state<=11;
					out<=238;
				end
				if(in == 837) begin
					state<=11;
					out<=239;
				end
				if(in == 838) begin
					state<=11;
					out<=240;
				end
				if(in == 839) begin
					state<=11;
					out<=241;
				end
				if(in == 840) begin
					state<=11;
					out<=242;
				end
				if(in == 841) begin
					state<=11;
					out<=243;
				end
				if(in == 842) begin
					state<=11;
					out<=244;
				end
				if(in == 843) begin
					state<=11;
					out<=245;
				end
				if(in == 844) begin
					state<=11;
					out<=246;
				end
				if(in == 845) begin
					state<=11;
					out<=247;
				end
				if(in == 846) begin
					state<=11;
					out<=248;
				end
				if(in == 847) begin
					state<=11;
					out<=249;
				end
				if(in == 848) begin
					state<=11;
					out<=250;
				end
				if(in == 849) begin
					state<=11;
					out<=251;
				end
				if(in == 850) begin
					state<=11;
					out<=252;
				end
				if(in == 851) begin
					state<=11;
					out<=253;
				end
				if(in == 852) begin
					state<=11;
					out<=254;
				end
				if(in == 853) begin
					state<=11;
					out<=255;
				end
				if(in == 854) begin
					state<=11;
					out<=0;
				end
				if(in == 855) begin
					state<=11;
					out<=1;
				end
				if(in == 856) begin
					state<=11;
					out<=2;
				end
				if(in == 857) begin
					state<=11;
					out<=3;
				end
				if(in == 858) begin
					state<=11;
					out<=4;
				end
				if(in == 859) begin
					state<=11;
					out<=5;
				end
				if(in == 860) begin
					state<=11;
					out<=6;
				end
				if(in == 861) begin
					state<=11;
					out<=7;
				end
				if(in == 862) begin
					state<=11;
					out<=8;
				end
				if(in == 863) begin
					state<=11;
					out<=9;
				end
				if(in == 864) begin
					state<=11;
					out<=10;
				end
				if(in == 865) begin
					state<=3;
					out<=11;
				end
				if(in == 866) begin
					state<=10;
					out<=12;
				end
				if(in == 867) begin
					state<=3;
					out<=13;
				end
				if(in == 868) begin
					state<=11;
					out<=14;
				end
				if(in == 869) begin
					state<=3;
					out<=15;
				end
				if(in == 870) begin
					state<=11;
					out<=16;
				end
				if(in == 871) begin
					state<=11;
					out<=17;
				end
				if(in == 872) begin
					state<=11;
					out<=18;
				end
				if(in == 873) begin
					state<=11;
					out<=19;
				end
				if(in == 874) begin
					state<=11;
					out<=20;
				end
				if(in == 875) begin
					state<=11;
					out<=21;
				end
				if(in == 876) begin
					state<=11;
					out<=22;
				end
				if(in == 877) begin
					state<=11;
					out<=23;
				end
				if(in == 878) begin
					state<=11;
					out<=24;
				end
				if(in == 879) begin
					state<=11;
					out<=25;
				end
				if(in == 880) begin
					state<=11;
					out<=26;
				end
				if(in == 881) begin
					state<=11;
					out<=27;
				end
				if(in == 882) begin
					state<=11;
					out<=28;
				end
				if(in == 883) begin
					state<=11;
					out<=29;
				end
				if(in == 884) begin
					state<=11;
					out<=30;
				end
				if(in == 885) begin
					state<=11;
					out<=31;
				end
				if(in == 886) begin
					state<=11;
					out<=32;
				end
				if(in == 887) begin
					state<=11;
					out<=33;
				end
				if(in == 888) begin
					state<=11;
					out<=34;
				end
				if(in == 889) begin
					state<=11;
					out<=35;
				end
				if(in == 890) begin
					state<=11;
					out<=36;
				end
				if(in == 891) begin
					state<=11;
					out<=37;
				end
				if(in == 892) begin
					state<=11;
					out<=38;
				end
				if(in == 893) begin
					state<=11;
					out<=39;
				end
				if(in == 894) begin
					state<=11;
					out<=40;
				end
				if(in == 895) begin
					state<=11;
					out<=41;
				end
				if(in == 896) begin
					state<=11;
					out<=42;
				end
				if(in == 897) begin
					state<=11;
					out<=43;
				end
				if(in == 898) begin
					state<=11;
					out<=44;
				end
				if(in == 899) begin
					state<=11;
					out<=45;
				end
				if(in == 900) begin
					state<=11;
					out<=46;
				end
				if(in == 901) begin
					state<=11;
					out<=47;
				end
				if(in == 902) begin
					state<=11;
					out<=48;
				end
				if(in == 903) begin
					state<=11;
					out<=49;
				end
				if(in == 904) begin
					state<=11;
					out<=50;
				end
				if(in == 905) begin
					state<=11;
					out<=51;
				end
				if(in == 906) begin
					state<=11;
					out<=52;
				end
				if(in == 907) begin
					state<=11;
					out<=53;
				end
				if(in == 908) begin
					state<=11;
					out<=54;
				end
				if(in == 909) begin
					state<=11;
					out<=55;
				end
				if(in == 910) begin
					state<=11;
					out<=56;
				end
				if(in == 911) begin
					state<=11;
					out<=57;
				end
				if(in == 912) begin
					state<=11;
					out<=58;
				end
				if(in == 913) begin
					state<=11;
					out<=59;
				end
				if(in == 914) begin
					state<=11;
					out<=60;
				end
				if(in == 915) begin
					state<=11;
					out<=61;
				end
				if(in == 916) begin
					state<=11;
					out<=62;
				end
				if(in == 917) begin
					state<=2;
					out<=63;
				end
				if(in == 918) begin
					state<=2;
					out<=64;
				end
				if(in == 919) begin
					state<=2;
					out<=65;
				end
				if(in == 920) begin
					state<=2;
					out<=66;
				end
				if(in == 921) begin
					state<=2;
					out<=67;
				end
				if(in == 922) begin
					state<=2;
					out<=68;
				end
				if(in == 923) begin
					state<=2;
					out<=69;
				end
				if(in == 924) begin
					state<=2;
					out<=70;
				end
				if(in == 925) begin
					state<=2;
					out<=71;
				end
				if(in == 926) begin
					state<=2;
					out<=72;
				end
				if(in == 927) begin
					state<=2;
					out<=73;
				end
				if(in == 928) begin
					state<=2;
					out<=74;
				end
			end
			11: begin
				if(in == 0) begin
					state<=3;
					out<=75;
				end
				if(in == 1) begin
					state<=1;
					out<=76;
				end
				if(in == 2) begin
					state<=11;
					out<=77;
				end
				if(in == 3) begin
					state<=3;
					out<=78;
				end
				if(in == 4) begin
					state<=12;
					out<=79;
				end
				if(in == 5) begin
					state<=3;
					out<=80;
				end
				if(in == 6) begin
					state<=12;
					out<=81;
				end
				if(in == 7) begin
					state<=12;
					out<=82;
				end
				if(in == 8) begin
					state<=12;
					out<=83;
				end
				if(in == 9) begin
					state<=12;
					out<=84;
				end
				if(in == 10) begin
					state<=12;
					out<=85;
				end
				if(in == 11) begin
					state<=12;
					out<=86;
				end
				if(in == 12) begin
					state<=12;
					out<=87;
				end
				if(in == 13) begin
					state<=12;
					out<=88;
				end
				if(in == 14) begin
					state<=12;
					out<=89;
				end
				if(in == 15) begin
					state<=12;
					out<=90;
				end
				if(in == 16) begin
					state<=12;
					out<=91;
				end
				if(in == 17) begin
					state<=12;
					out<=92;
				end
				if(in == 18) begin
					state<=12;
					out<=93;
				end
				if(in == 19) begin
					state<=12;
					out<=94;
				end
				if(in == 20) begin
					state<=12;
					out<=95;
				end
				if(in == 21) begin
					state<=12;
					out<=96;
				end
				if(in == 22) begin
					state<=12;
					out<=97;
				end
				if(in == 23) begin
					state<=12;
					out<=98;
				end
				if(in == 24) begin
					state<=12;
					out<=99;
				end
				if(in == 25) begin
					state<=12;
					out<=100;
				end
				if(in == 26) begin
					state<=12;
					out<=101;
				end
				if(in == 27) begin
					state<=12;
					out<=102;
				end
				if(in == 28) begin
					state<=12;
					out<=103;
				end
				if(in == 29) begin
					state<=12;
					out<=104;
				end
				if(in == 30) begin
					state<=12;
					out<=105;
				end
				if(in == 31) begin
					state<=12;
					out<=106;
				end
				if(in == 32) begin
					state<=12;
					out<=107;
				end
				if(in == 33) begin
					state<=12;
					out<=108;
				end
				if(in == 34) begin
					state<=12;
					out<=109;
				end
				if(in == 35) begin
					state<=12;
					out<=110;
				end
				if(in == 36) begin
					state<=12;
					out<=111;
				end
				if(in == 37) begin
					state<=12;
					out<=112;
				end
				if(in == 38) begin
					state<=12;
					out<=113;
				end
				if(in == 39) begin
					state<=12;
					out<=114;
				end
				if(in == 40) begin
					state<=12;
					out<=115;
				end
				if(in == 41) begin
					state<=12;
					out<=116;
				end
				if(in == 42) begin
					state<=12;
					out<=117;
				end
				if(in == 43) begin
					state<=12;
					out<=118;
				end
				if(in == 44) begin
					state<=12;
					out<=119;
				end
				if(in == 45) begin
					state<=12;
					out<=120;
				end
				if(in == 46) begin
					state<=12;
					out<=121;
				end
				if(in == 47) begin
					state<=12;
					out<=122;
				end
				if(in == 48) begin
					state<=12;
					out<=123;
				end
				if(in == 49) begin
					state<=12;
					out<=124;
				end
				if(in == 50) begin
					state<=12;
					out<=125;
				end
				if(in == 51) begin
					state<=12;
					out<=126;
				end
				if(in == 52) begin
					state<=12;
					out<=127;
				end
				if(in == 53) begin
					state<=3;
					out<=128;
				end
				if(in == 54) begin
					state<=11;
					out<=129;
				end
				if(in == 55) begin
					state<=3;
					out<=130;
				end
				if(in == 56) begin
					state<=12;
					out<=131;
				end
				if(in == 57) begin
					state<=3;
					out<=132;
				end
				if(in == 58) begin
					state<=12;
					out<=133;
				end
				if(in == 59) begin
					state<=12;
					out<=134;
				end
				if(in == 60) begin
					state<=12;
					out<=135;
				end
				if(in == 61) begin
					state<=12;
					out<=136;
				end
				if(in == 62) begin
					state<=12;
					out<=137;
				end
				if(in == 63) begin
					state<=12;
					out<=138;
				end
				if(in == 64) begin
					state<=12;
					out<=139;
				end
				if(in == 65) begin
					state<=12;
					out<=140;
				end
				if(in == 66) begin
					state<=12;
					out<=141;
				end
				if(in == 67) begin
					state<=12;
					out<=142;
				end
				if(in == 68) begin
					state<=12;
					out<=143;
				end
				if(in == 69) begin
					state<=12;
					out<=144;
				end
				if(in == 70) begin
					state<=12;
					out<=145;
				end
				if(in == 71) begin
					state<=12;
					out<=146;
				end
				if(in == 72) begin
					state<=12;
					out<=147;
				end
				if(in == 73) begin
					state<=12;
					out<=148;
				end
				if(in == 74) begin
					state<=12;
					out<=149;
				end
				if(in == 75) begin
					state<=12;
					out<=150;
				end
				if(in == 76) begin
					state<=12;
					out<=151;
				end
				if(in == 77) begin
					state<=12;
					out<=152;
				end
				if(in == 78) begin
					state<=12;
					out<=153;
				end
				if(in == 79) begin
					state<=12;
					out<=154;
				end
				if(in == 80) begin
					state<=12;
					out<=155;
				end
				if(in == 81) begin
					state<=12;
					out<=156;
				end
				if(in == 82) begin
					state<=12;
					out<=157;
				end
				if(in == 83) begin
					state<=12;
					out<=158;
				end
				if(in == 84) begin
					state<=12;
					out<=159;
				end
				if(in == 85) begin
					state<=12;
					out<=160;
				end
				if(in == 86) begin
					state<=12;
					out<=161;
				end
				if(in == 87) begin
					state<=12;
					out<=162;
				end
				if(in == 88) begin
					state<=12;
					out<=163;
				end
				if(in == 89) begin
					state<=12;
					out<=164;
				end
				if(in == 90) begin
					state<=12;
					out<=165;
				end
				if(in == 91) begin
					state<=12;
					out<=166;
				end
				if(in == 92) begin
					state<=12;
					out<=167;
				end
				if(in == 93) begin
					state<=12;
					out<=168;
				end
				if(in == 94) begin
					state<=12;
					out<=169;
				end
				if(in == 95) begin
					state<=12;
					out<=170;
				end
				if(in == 96) begin
					state<=12;
					out<=171;
				end
				if(in == 97) begin
					state<=12;
					out<=172;
				end
				if(in == 98) begin
					state<=12;
					out<=173;
				end
				if(in == 99) begin
					state<=12;
					out<=174;
				end
				if(in == 100) begin
					state<=12;
					out<=175;
				end
				if(in == 101) begin
					state<=12;
					out<=176;
				end
				if(in == 102) begin
					state<=12;
					out<=177;
				end
				if(in == 103) begin
					state<=12;
					out<=178;
				end
				if(in == 104) begin
					state<=12;
					out<=179;
				end
				if(in == 105) begin
					state<=2;
					out<=180;
				end
				if(in == 106) begin
					state<=2;
					out<=181;
				end
				if(in == 107) begin
					state<=2;
					out<=182;
				end
				if(in == 108) begin
					state<=2;
					out<=183;
				end
				if(in == 109) begin
					state<=2;
					out<=184;
				end
				if(in == 110) begin
					state<=2;
					out<=185;
				end
				if(in == 111) begin
					state<=2;
					out<=186;
				end
				if(in == 112) begin
					state<=2;
					out<=187;
				end
				if(in == 113) begin
					state<=2;
					out<=188;
				end
				if(in == 114) begin
					state<=2;
					out<=189;
				end
				if(in == 115) begin
					state<=2;
					out<=190;
				end
				if(in == 116) begin
					state<=2;
					out<=191;
				end
				if(in == 117) begin
					state<=3;
					out<=192;
				end
				if(in == 118) begin
					state<=11;
					out<=193;
				end
				if(in == 119) begin
					state<=3;
					out<=194;
				end
				if(in == 120) begin
					state<=12;
					out<=195;
				end
				if(in == 121) begin
					state<=3;
					out<=196;
				end
				if(in == 122) begin
					state<=12;
					out<=197;
				end
				if(in == 123) begin
					state<=12;
					out<=198;
				end
				if(in == 124) begin
					state<=12;
					out<=199;
				end
				if(in == 125) begin
					state<=12;
					out<=200;
				end
				if(in == 126) begin
					state<=12;
					out<=201;
				end
				if(in == 127) begin
					state<=12;
					out<=202;
				end
				if(in == 128) begin
					state<=12;
					out<=203;
				end
				if(in == 129) begin
					state<=12;
					out<=204;
				end
				if(in == 130) begin
					state<=12;
					out<=205;
				end
				if(in == 131) begin
					state<=12;
					out<=206;
				end
				if(in == 132) begin
					state<=12;
					out<=207;
				end
				if(in == 133) begin
					state<=12;
					out<=208;
				end
				if(in == 134) begin
					state<=12;
					out<=209;
				end
				if(in == 135) begin
					state<=12;
					out<=210;
				end
				if(in == 136) begin
					state<=12;
					out<=211;
				end
				if(in == 137) begin
					state<=12;
					out<=212;
				end
				if(in == 138) begin
					state<=12;
					out<=213;
				end
				if(in == 139) begin
					state<=12;
					out<=214;
				end
				if(in == 140) begin
					state<=12;
					out<=215;
				end
				if(in == 141) begin
					state<=12;
					out<=216;
				end
				if(in == 142) begin
					state<=12;
					out<=217;
				end
				if(in == 143) begin
					state<=12;
					out<=218;
				end
				if(in == 144) begin
					state<=12;
					out<=219;
				end
				if(in == 145) begin
					state<=12;
					out<=220;
				end
				if(in == 146) begin
					state<=12;
					out<=221;
				end
				if(in == 147) begin
					state<=12;
					out<=222;
				end
				if(in == 148) begin
					state<=12;
					out<=223;
				end
				if(in == 149) begin
					state<=12;
					out<=224;
				end
				if(in == 150) begin
					state<=12;
					out<=225;
				end
				if(in == 151) begin
					state<=12;
					out<=226;
				end
				if(in == 152) begin
					state<=12;
					out<=227;
				end
				if(in == 153) begin
					state<=12;
					out<=228;
				end
				if(in == 154) begin
					state<=12;
					out<=229;
				end
				if(in == 155) begin
					state<=12;
					out<=230;
				end
				if(in == 156) begin
					state<=12;
					out<=231;
				end
				if(in == 157) begin
					state<=12;
					out<=232;
				end
				if(in == 158) begin
					state<=12;
					out<=233;
				end
				if(in == 159) begin
					state<=12;
					out<=234;
				end
				if(in == 160) begin
					state<=12;
					out<=235;
				end
				if(in == 161) begin
					state<=12;
					out<=236;
				end
				if(in == 162) begin
					state<=12;
					out<=237;
				end
				if(in == 163) begin
					state<=12;
					out<=238;
				end
				if(in == 164) begin
					state<=12;
					out<=239;
				end
				if(in == 165) begin
					state<=12;
					out<=240;
				end
				if(in == 166) begin
					state<=12;
					out<=241;
				end
				if(in == 167) begin
					state<=12;
					out<=242;
				end
				if(in == 168) begin
					state<=12;
					out<=243;
				end
				if(in == 169) begin
					state<=3;
					out<=244;
				end
				if(in == 170) begin
					state<=11;
					out<=245;
				end
				if(in == 171) begin
					state<=3;
					out<=246;
				end
				if(in == 172) begin
					state<=12;
					out<=247;
				end
				if(in == 173) begin
					state<=3;
					out<=248;
				end
				if(in == 174) begin
					state<=12;
					out<=249;
				end
				if(in == 175) begin
					state<=12;
					out<=250;
				end
				if(in == 176) begin
					state<=12;
					out<=251;
				end
				if(in == 177) begin
					state<=12;
					out<=252;
				end
				if(in == 178) begin
					state<=12;
					out<=253;
				end
				if(in == 179) begin
					state<=12;
					out<=254;
				end
				if(in == 180) begin
					state<=12;
					out<=255;
				end
				if(in == 181) begin
					state<=12;
					out<=0;
				end
				if(in == 182) begin
					state<=12;
					out<=1;
				end
				if(in == 183) begin
					state<=12;
					out<=2;
				end
				if(in == 184) begin
					state<=12;
					out<=3;
				end
				if(in == 185) begin
					state<=12;
					out<=4;
				end
				if(in == 186) begin
					state<=12;
					out<=5;
				end
				if(in == 187) begin
					state<=12;
					out<=6;
				end
				if(in == 188) begin
					state<=12;
					out<=7;
				end
				if(in == 189) begin
					state<=12;
					out<=8;
				end
				if(in == 190) begin
					state<=12;
					out<=9;
				end
				if(in == 191) begin
					state<=12;
					out<=10;
				end
				if(in == 192) begin
					state<=12;
					out<=11;
				end
				if(in == 193) begin
					state<=12;
					out<=12;
				end
				if(in == 194) begin
					state<=12;
					out<=13;
				end
				if(in == 195) begin
					state<=12;
					out<=14;
				end
				if(in == 196) begin
					state<=12;
					out<=15;
				end
				if(in == 197) begin
					state<=12;
					out<=16;
				end
				if(in == 198) begin
					state<=12;
					out<=17;
				end
				if(in == 199) begin
					state<=12;
					out<=18;
				end
				if(in == 200) begin
					state<=12;
					out<=19;
				end
				if(in == 201) begin
					state<=12;
					out<=20;
				end
				if(in == 202) begin
					state<=12;
					out<=21;
				end
				if(in == 203) begin
					state<=12;
					out<=22;
				end
				if(in == 204) begin
					state<=12;
					out<=23;
				end
				if(in == 205) begin
					state<=12;
					out<=24;
				end
				if(in == 206) begin
					state<=12;
					out<=25;
				end
				if(in == 207) begin
					state<=12;
					out<=26;
				end
				if(in == 208) begin
					state<=12;
					out<=27;
				end
				if(in == 209) begin
					state<=12;
					out<=28;
				end
				if(in == 210) begin
					state<=12;
					out<=29;
				end
				if(in == 211) begin
					state<=12;
					out<=30;
				end
				if(in == 212) begin
					state<=12;
					out<=31;
				end
				if(in == 213) begin
					state<=12;
					out<=32;
				end
				if(in == 214) begin
					state<=12;
					out<=33;
				end
				if(in == 215) begin
					state<=12;
					out<=34;
				end
				if(in == 216) begin
					state<=12;
					out<=35;
				end
				if(in == 217) begin
					state<=12;
					out<=36;
				end
				if(in == 218) begin
					state<=12;
					out<=37;
				end
				if(in == 219) begin
					state<=12;
					out<=38;
				end
				if(in == 220) begin
					state<=12;
					out<=39;
				end
				if(in == 221) begin
					state<=2;
					out<=40;
				end
				if(in == 222) begin
					state<=2;
					out<=41;
				end
				if(in == 223) begin
					state<=2;
					out<=42;
				end
				if(in == 224) begin
					state<=2;
					out<=43;
				end
				if(in == 225) begin
					state<=2;
					out<=44;
				end
				if(in == 226) begin
					state<=2;
					out<=45;
				end
				if(in == 227) begin
					state<=2;
					out<=46;
				end
				if(in == 228) begin
					state<=2;
					out<=47;
				end
				if(in == 229) begin
					state<=2;
					out<=48;
				end
				if(in == 230) begin
					state<=2;
					out<=49;
				end
				if(in == 231) begin
					state<=2;
					out<=50;
				end
				if(in == 232) begin
					state<=2;
					out<=51;
				end
				if(in == 233) begin
					state<=3;
					out<=52;
				end
				if(in == 234) begin
					state<=11;
					out<=53;
				end
				if(in == 235) begin
					state<=3;
					out<=54;
				end
				if(in == 236) begin
					state<=12;
					out<=55;
				end
				if(in == 237) begin
					state<=3;
					out<=56;
				end
				if(in == 238) begin
					state<=12;
					out<=57;
				end
				if(in == 239) begin
					state<=12;
					out<=58;
				end
				if(in == 240) begin
					state<=12;
					out<=59;
				end
				if(in == 241) begin
					state<=12;
					out<=60;
				end
				if(in == 242) begin
					state<=12;
					out<=61;
				end
				if(in == 243) begin
					state<=12;
					out<=62;
				end
				if(in == 244) begin
					state<=12;
					out<=63;
				end
				if(in == 245) begin
					state<=12;
					out<=64;
				end
				if(in == 246) begin
					state<=12;
					out<=65;
				end
				if(in == 247) begin
					state<=12;
					out<=66;
				end
				if(in == 248) begin
					state<=12;
					out<=67;
				end
				if(in == 249) begin
					state<=12;
					out<=68;
				end
				if(in == 250) begin
					state<=12;
					out<=69;
				end
				if(in == 251) begin
					state<=12;
					out<=70;
				end
				if(in == 252) begin
					state<=12;
					out<=71;
				end
				if(in == 253) begin
					state<=12;
					out<=72;
				end
				if(in == 254) begin
					state<=12;
					out<=73;
				end
				if(in == 255) begin
					state<=12;
					out<=74;
				end
				if(in == 256) begin
					state<=12;
					out<=75;
				end
				if(in == 257) begin
					state<=12;
					out<=76;
				end
				if(in == 258) begin
					state<=12;
					out<=77;
				end
				if(in == 259) begin
					state<=12;
					out<=78;
				end
				if(in == 260) begin
					state<=12;
					out<=79;
				end
				if(in == 261) begin
					state<=12;
					out<=80;
				end
				if(in == 262) begin
					state<=12;
					out<=81;
				end
				if(in == 263) begin
					state<=12;
					out<=82;
				end
				if(in == 264) begin
					state<=12;
					out<=83;
				end
				if(in == 265) begin
					state<=12;
					out<=84;
				end
				if(in == 266) begin
					state<=12;
					out<=85;
				end
				if(in == 267) begin
					state<=12;
					out<=86;
				end
				if(in == 268) begin
					state<=12;
					out<=87;
				end
				if(in == 269) begin
					state<=12;
					out<=88;
				end
				if(in == 270) begin
					state<=12;
					out<=89;
				end
				if(in == 271) begin
					state<=12;
					out<=90;
				end
				if(in == 272) begin
					state<=12;
					out<=91;
				end
				if(in == 273) begin
					state<=12;
					out<=92;
				end
				if(in == 274) begin
					state<=12;
					out<=93;
				end
				if(in == 275) begin
					state<=12;
					out<=94;
				end
				if(in == 276) begin
					state<=12;
					out<=95;
				end
				if(in == 277) begin
					state<=12;
					out<=96;
				end
				if(in == 278) begin
					state<=12;
					out<=97;
				end
				if(in == 279) begin
					state<=12;
					out<=98;
				end
				if(in == 280) begin
					state<=12;
					out<=99;
				end
				if(in == 281) begin
					state<=12;
					out<=100;
				end
				if(in == 282) begin
					state<=12;
					out<=101;
				end
				if(in == 283) begin
					state<=12;
					out<=102;
				end
				if(in == 284) begin
					state<=12;
					out<=103;
				end
				if(in == 285) begin
					state<=3;
					out<=104;
				end
				if(in == 286) begin
					state<=11;
					out<=105;
				end
				if(in == 287) begin
					state<=3;
					out<=106;
				end
				if(in == 288) begin
					state<=12;
					out<=107;
				end
				if(in == 289) begin
					state<=3;
					out<=108;
				end
				if(in == 290) begin
					state<=12;
					out<=109;
				end
				if(in == 291) begin
					state<=12;
					out<=110;
				end
				if(in == 292) begin
					state<=12;
					out<=111;
				end
				if(in == 293) begin
					state<=12;
					out<=112;
				end
				if(in == 294) begin
					state<=12;
					out<=113;
				end
				if(in == 295) begin
					state<=12;
					out<=114;
				end
				if(in == 296) begin
					state<=12;
					out<=115;
				end
				if(in == 297) begin
					state<=12;
					out<=116;
				end
				if(in == 298) begin
					state<=12;
					out<=117;
				end
				if(in == 299) begin
					state<=12;
					out<=118;
				end
				if(in == 300) begin
					state<=12;
					out<=119;
				end
				if(in == 301) begin
					state<=12;
					out<=120;
				end
				if(in == 302) begin
					state<=12;
					out<=121;
				end
				if(in == 303) begin
					state<=12;
					out<=122;
				end
				if(in == 304) begin
					state<=12;
					out<=123;
				end
				if(in == 305) begin
					state<=12;
					out<=124;
				end
				if(in == 306) begin
					state<=12;
					out<=125;
				end
				if(in == 307) begin
					state<=12;
					out<=126;
				end
				if(in == 308) begin
					state<=12;
					out<=127;
				end
				if(in == 309) begin
					state<=12;
					out<=128;
				end
				if(in == 310) begin
					state<=12;
					out<=129;
				end
				if(in == 311) begin
					state<=12;
					out<=130;
				end
				if(in == 312) begin
					state<=12;
					out<=131;
				end
				if(in == 313) begin
					state<=12;
					out<=132;
				end
				if(in == 314) begin
					state<=12;
					out<=133;
				end
				if(in == 315) begin
					state<=12;
					out<=134;
				end
				if(in == 316) begin
					state<=12;
					out<=135;
				end
				if(in == 317) begin
					state<=12;
					out<=136;
				end
				if(in == 318) begin
					state<=12;
					out<=137;
				end
				if(in == 319) begin
					state<=12;
					out<=138;
				end
				if(in == 320) begin
					state<=12;
					out<=139;
				end
				if(in == 321) begin
					state<=12;
					out<=140;
				end
				if(in == 322) begin
					state<=12;
					out<=141;
				end
				if(in == 323) begin
					state<=12;
					out<=142;
				end
				if(in == 324) begin
					state<=12;
					out<=143;
				end
				if(in == 325) begin
					state<=12;
					out<=144;
				end
				if(in == 326) begin
					state<=12;
					out<=145;
				end
				if(in == 327) begin
					state<=12;
					out<=146;
				end
				if(in == 328) begin
					state<=12;
					out<=147;
				end
				if(in == 329) begin
					state<=12;
					out<=148;
				end
				if(in == 330) begin
					state<=12;
					out<=149;
				end
				if(in == 331) begin
					state<=12;
					out<=150;
				end
				if(in == 332) begin
					state<=12;
					out<=151;
				end
				if(in == 333) begin
					state<=12;
					out<=152;
				end
				if(in == 334) begin
					state<=12;
					out<=153;
				end
				if(in == 335) begin
					state<=12;
					out<=154;
				end
				if(in == 336) begin
					state<=12;
					out<=155;
				end
				if(in == 337) begin
					state<=2;
					out<=156;
				end
				if(in == 338) begin
					state<=2;
					out<=157;
				end
				if(in == 339) begin
					state<=2;
					out<=158;
				end
				if(in == 340) begin
					state<=2;
					out<=159;
				end
				if(in == 341) begin
					state<=2;
					out<=160;
				end
				if(in == 342) begin
					state<=2;
					out<=161;
				end
				if(in == 343) begin
					state<=2;
					out<=162;
				end
				if(in == 344) begin
					state<=2;
					out<=163;
				end
				if(in == 345) begin
					state<=2;
					out<=164;
				end
				if(in == 346) begin
					state<=2;
					out<=165;
				end
				if(in == 347) begin
					state<=2;
					out<=166;
				end
				if(in == 348) begin
					state<=2;
					out<=167;
				end
				if(in == 349) begin
					state<=3;
					out<=168;
				end
				if(in == 350) begin
					state<=11;
					out<=169;
				end
				if(in == 351) begin
					state<=3;
					out<=170;
				end
				if(in == 352) begin
					state<=12;
					out<=171;
				end
				if(in == 353) begin
					state<=3;
					out<=172;
				end
				if(in == 354) begin
					state<=12;
					out<=173;
				end
				if(in == 355) begin
					state<=12;
					out<=174;
				end
				if(in == 356) begin
					state<=12;
					out<=175;
				end
				if(in == 357) begin
					state<=12;
					out<=176;
				end
				if(in == 358) begin
					state<=12;
					out<=177;
				end
				if(in == 359) begin
					state<=12;
					out<=178;
				end
				if(in == 360) begin
					state<=12;
					out<=179;
				end
				if(in == 361) begin
					state<=12;
					out<=180;
				end
				if(in == 362) begin
					state<=12;
					out<=181;
				end
				if(in == 363) begin
					state<=12;
					out<=182;
				end
				if(in == 364) begin
					state<=12;
					out<=183;
				end
				if(in == 365) begin
					state<=12;
					out<=184;
				end
				if(in == 366) begin
					state<=12;
					out<=185;
				end
				if(in == 367) begin
					state<=12;
					out<=186;
				end
				if(in == 368) begin
					state<=12;
					out<=187;
				end
				if(in == 369) begin
					state<=12;
					out<=188;
				end
				if(in == 370) begin
					state<=12;
					out<=189;
				end
				if(in == 371) begin
					state<=12;
					out<=190;
				end
				if(in == 372) begin
					state<=12;
					out<=191;
				end
				if(in == 373) begin
					state<=12;
					out<=192;
				end
				if(in == 374) begin
					state<=12;
					out<=193;
				end
				if(in == 375) begin
					state<=12;
					out<=194;
				end
				if(in == 376) begin
					state<=12;
					out<=195;
				end
				if(in == 377) begin
					state<=12;
					out<=196;
				end
				if(in == 378) begin
					state<=12;
					out<=197;
				end
				if(in == 379) begin
					state<=12;
					out<=198;
				end
				if(in == 380) begin
					state<=12;
					out<=199;
				end
				if(in == 381) begin
					state<=12;
					out<=200;
				end
				if(in == 382) begin
					state<=12;
					out<=201;
				end
				if(in == 383) begin
					state<=12;
					out<=202;
				end
				if(in == 384) begin
					state<=12;
					out<=203;
				end
				if(in == 385) begin
					state<=12;
					out<=204;
				end
				if(in == 386) begin
					state<=12;
					out<=205;
				end
				if(in == 387) begin
					state<=12;
					out<=206;
				end
				if(in == 388) begin
					state<=12;
					out<=207;
				end
				if(in == 389) begin
					state<=12;
					out<=208;
				end
				if(in == 390) begin
					state<=12;
					out<=209;
				end
				if(in == 391) begin
					state<=12;
					out<=210;
				end
				if(in == 392) begin
					state<=12;
					out<=211;
				end
				if(in == 393) begin
					state<=12;
					out<=212;
				end
				if(in == 394) begin
					state<=12;
					out<=213;
				end
				if(in == 395) begin
					state<=12;
					out<=214;
				end
				if(in == 396) begin
					state<=12;
					out<=215;
				end
				if(in == 397) begin
					state<=12;
					out<=216;
				end
				if(in == 398) begin
					state<=12;
					out<=217;
				end
				if(in == 399) begin
					state<=12;
					out<=218;
				end
				if(in == 400) begin
					state<=12;
					out<=219;
				end
				if(in == 401) begin
					state<=3;
					out<=220;
				end
				if(in == 402) begin
					state<=11;
					out<=221;
				end
				if(in == 403) begin
					state<=3;
					out<=222;
				end
				if(in == 404) begin
					state<=12;
					out<=223;
				end
				if(in == 405) begin
					state<=3;
					out<=224;
				end
				if(in == 406) begin
					state<=12;
					out<=225;
				end
				if(in == 407) begin
					state<=12;
					out<=226;
				end
				if(in == 408) begin
					state<=12;
					out<=227;
				end
				if(in == 409) begin
					state<=12;
					out<=228;
				end
				if(in == 410) begin
					state<=12;
					out<=229;
				end
				if(in == 411) begin
					state<=12;
					out<=230;
				end
				if(in == 412) begin
					state<=12;
					out<=231;
				end
				if(in == 413) begin
					state<=12;
					out<=232;
				end
				if(in == 414) begin
					state<=12;
					out<=233;
				end
				if(in == 415) begin
					state<=12;
					out<=234;
				end
				if(in == 416) begin
					state<=12;
					out<=235;
				end
				if(in == 417) begin
					state<=12;
					out<=236;
				end
				if(in == 418) begin
					state<=12;
					out<=237;
				end
				if(in == 419) begin
					state<=12;
					out<=238;
				end
				if(in == 420) begin
					state<=12;
					out<=239;
				end
				if(in == 421) begin
					state<=12;
					out<=240;
				end
				if(in == 422) begin
					state<=12;
					out<=241;
				end
				if(in == 423) begin
					state<=12;
					out<=242;
				end
				if(in == 424) begin
					state<=12;
					out<=243;
				end
				if(in == 425) begin
					state<=12;
					out<=244;
				end
				if(in == 426) begin
					state<=12;
					out<=245;
				end
				if(in == 427) begin
					state<=12;
					out<=246;
				end
				if(in == 428) begin
					state<=12;
					out<=247;
				end
				if(in == 429) begin
					state<=12;
					out<=248;
				end
				if(in == 430) begin
					state<=12;
					out<=249;
				end
				if(in == 431) begin
					state<=12;
					out<=250;
				end
				if(in == 432) begin
					state<=12;
					out<=251;
				end
				if(in == 433) begin
					state<=12;
					out<=252;
				end
				if(in == 434) begin
					state<=12;
					out<=253;
				end
				if(in == 435) begin
					state<=12;
					out<=254;
				end
				if(in == 436) begin
					state<=12;
					out<=255;
				end
				if(in == 437) begin
					state<=12;
					out<=0;
				end
				if(in == 438) begin
					state<=12;
					out<=1;
				end
				if(in == 439) begin
					state<=12;
					out<=2;
				end
				if(in == 440) begin
					state<=12;
					out<=3;
				end
				if(in == 441) begin
					state<=12;
					out<=4;
				end
				if(in == 442) begin
					state<=12;
					out<=5;
				end
				if(in == 443) begin
					state<=12;
					out<=6;
				end
				if(in == 444) begin
					state<=12;
					out<=7;
				end
				if(in == 445) begin
					state<=12;
					out<=8;
				end
				if(in == 446) begin
					state<=12;
					out<=9;
				end
				if(in == 447) begin
					state<=12;
					out<=10;
				end
				if(in == 448) begin
					state<=12;
					out<=11;
				end
				if(in == 449) begin
					state<=12;
					out<=12;
				end
				if(in == 450) begin
					state<=12;
					out<=13;
				end
				if(in == 451) begin
					state<=12;
					out<=14;
				end
				if(in == 452) begin
					state<=12;
					out<=15;
				end
				if(in == 453) begin
					state<=2;
					out<=16;
				end
				if(in == 454) begin
					state<=2;
					out<=17;
				end
				if(in == 455) begin
					state<=2;
					out<=18;
				end
				if(in == 456) begin
					state<=2;
					out<=19;
				end
				if(in == 457) begin
					state<=2;
					out<=20;
				end
				if(in == 458) begin
					state<=2;
					out<=21;
				end
				if(in == 459) begin
					state<=2;
					out<=22;
				end
				if(in == 460) begin
					state<=2;
					out<=23;
				end
				if(in == 461) begin
					state<=2;
					out<=24;
				end
				if(in == 462) begin
					state<=2;
					out<=25;
				end
				if(in == 463) begin
					state<=2;
					out<=26;
				end
				if(in == 464) begin
					state<=2;
					out<=27;
				end
				if(in == 465) begin
					state<=3;
					out<=28;
				end
				if(in == 466) begin
					state<=11;
					out<=29;
				end
				if(in == 467) begin
					state<=3;
					out<=30;
				end
				if(in == 468) begin
					state<=12;
					out<=31;
				end
				if(in == 469) begin
					state<=3;
					out<=32;
				end
				if(in == 470) begin
					state<=12;
					out<=33;
				end
				if(in == 471) begin
					state<=12;
					out<=34;
				end
				if(in == 472) begin
					state<=12;
					out<=35;
				end
				if(in == 473) begin
					state<=12;
					out<=36;
				end
				if(in == 474) begin
					state<=12;
					out<=37;
				end
				if(in == 475) begin
					state<=12;
					out<=38;
				end
				if(in == 476) begin
					state<=12;
					out<=39;
				end
				if(in == 477) begin
					state<=12;
					out<=40;
				end
				if(in == 478) begin
					state<=12;
					out<=41;
				end
				if(in == 479) begin
					state<=12;
					out<=42;
				end
				if(in == 480) begin
					state<=12;
					out<=43;
				end
				if(in == 481) begin
					state<=12;
					out<=44;
				end
				if(in == 482) begin
					state<=12;
					out<=45;
				end
				if(in == 483) begin
					state<=12;
					out<=46;
				end
				if(in == 484) begin
					state<=12;
					out<=47;
				end
				if(in == 485) begin
					state<=12;
					out<=48;
				end
				if(in == 486) begin
					state<=12;
					out<=49;
				end
				if(in == 487) begin
					state<=12;
					out<=50;
				end
				if(in == 488) begin
					state<=12;
					out<=51;
				end
				if(in == 489) begin
					state<=12;
					out<=52;
				end
				if(in == 490) begin
					state<=12;
					out<=53;
				end
				if(in == 491) begin
					state<=12;
					out<=54;
				end
				if(in == 492) begin
					state<=12;
					out<=55;
				end
				if(in == 493) begin
					state<=12;
					out<=56;
				end
				if(in == 494) begin
					state<=12;
					out<=57;
				end
				if(in == 495) begin
					state<=12;
					out<=58;
				end
				if(in == 496) begin
					state<=12;
					out<=59;
				end
				if(in == 497) begin
					state<=12;
					out<=60;
				end
				if(in == 498) begin
					state<=12;
					out<=61;
				end
				if(in == 499) begin
					state<=12;
					out<=62;
				end
				if(in == 500) begin
					state<=12;
					out<=63;
				end
				if(in == 501) begin
					state<=12;
					out<=64;
				end
				if(in == 502) begin
					state<=12;
					out<=65;
				end
				if(in == 503) begin
					state<=12;
					out<=66;
				end
				if(in == 504) begin
					state<=12;
					out<=67;
				end
				if(in == 505) begin
					state<=12;
					out<=68;
				end
				if(in == 506) begin
					state<=12;
					out<=69;
				end
				if(in == 507) begin
					state<=12;
					out<=70;
				end
				if(in == 508) begin
					state<=12;
					out<=71;
				end
				if(in == 509) begin
					state<=12;
					out<=72;
				end
				if(in == 510) begin
					state<=12;
					out<=73;
				end
				if(in == 511) begin
					state<=12;
					out<=74;
				end
				if(in == 512) begin
					state<=12;
					out<=75;
				end
				if(in == 513) begin
					state<=12;
					out<=76;
				end
				if(in == 514) begin
					state<=12;
					out<=77;
				end
				if(in == 515) begin
					state<=12;
					out<=78;
				end
				if(in == 516) begin
					state<=12;
					out<=79;
				end
				if(in == 517) begin
					state<=3;
					out<=80;
				end
				if(in == 518) begin
					state<=11;
					out<=81;
				end
				if(in == 519) begin
					state<=3;
					out<=82;
				end
				if(in == 520) begin
					state<=12;
					out<=83;
				end
				if(in == 521) begin
					state<=3;
					out<=84;
				end
				if(in == 522) begin
					state<=12;
					out<=85;
				end
				if(in == 523) begin
					state<=12;
					out<=86;
				end
				if(in == 524) begin
					state<=12;
					out<=87;
				end
				if(in == 525) begin
					state<=12;
					out<=88;
				end
				if(in == 526) begin
					state<=12;
					out<=89;
				end
				if(in == 527) begin
					state<=12;
					out<=90;
				end
				if(in == 528) begin
					state<=12;
					out<=91;
				end
				if(in == 529) begin
					state<=12;
					out<=92;
				end
				if(in == 530) begin
					state<=12;
					out<=93;
				end
				if(in == 531) begin
					state<=12;
					out<=94;
				end
				if(in == 532) begin
					state<=12;
					out<=95;
				end
				if(in == 533) begin
					state<=12;
					out<=96;
				end
				if(in == 534) begin
					state<=12;
					out<=97;
				end
				if(in == 535) begin
					state<=12;
					out<=98;
				end
				if(in == 536) begin
					state<=12;
					out<=99;
				end
				if(in == 537) begin
					state<=12;
					out<=100;
				end
				if(in == 538) begin
					state<=12;
					out<=101;
				end
				if(in == 539) begin
					state<=12;
					out<=102;
				end
				if(in == 540) begin
					state<=12;
					out<=103;
				end
				if(in == 541) begin
					state<=12;
					out<=104;
				end
				if(in == 542) begin
					state<=12;
					out<=105;
				end
				if(in == 543) begin
					state<=12;
					out<=106;
				end
				if(in == 544) begin
					state<=12;
					out<=107;
				end
				if(in == 545) begin
					state<=12;
					out<=108;
				end
				if(in == 546) begin
					state<=12;
					out<=109;
				end
				if(in == 547) begin
					state<=12;
					out<=110;
				end
				if(in == 548) begin
					state<=12;
					out<=111;
				end
				if(in == 549) begin
					state<=12;
					out<=112;
				end
				if(in == 550) begin
					state<=12;
					out<=113;
				end
				if(in == 551) begin
					state<=12;
					out<=114;
				end
				if(in == 552) begin
					state<=12;
					out<=115;
				end
				if(in == 553) begin
					state<=12;
					out<=116;
				end
				if(in == 554) begin
					state<=12;
					out<=117;
				end
				if(in == 555) begin
					state<=12;
					out<=118;
				end
				if(in == 556) begin
					state<=12;
					out<=119;
				end
				if(in == 557) begin
					state<=12;
					out<=120;
				end
				if(in == 558) begin
					state<=12;
					out<=121;
				end
				if(in == 559) begin
					state<=12;
					out<=122;
				end
				if(in == 560) begin
					state<=12;
					out<=123;
				end
				if(in == 561) begin
					state<=12;
					out<=124;
				end
				if(in == 562) begin
					state<=12;
					out<=125;
				end
				if(in == 563) begin
					state<=12;
					out<=126;
				end
				if(in == 564) begin
					state<=12;
					out<=127;
				end
				if(in == 565) begin
					state<=12;
					out<=128;
				end
				if(in == 566) begin
					state<=12;
					out<=129;
				end
				if(in == 567) begin
					state<=12;
					out<=130;
				end
				if(in == 568) begin
					state<=12;
					out<=131;
				end
				if(in == 569) begin
					state<=2;
					out<=132;
				end
				if(in == 570) begin
					state<=2;
					out<=133;
				end
				if(in == 571) begin
					state<=2;
					out<=134;
				end
				if(in == 572) begin
					state<=2;
					out<=135;
				end
				if(in == 573) begin
					state<=2;
					out<=136;
				end
				if(in == 574) begin
					state<=2;
					out<=137;
				end
				if(in == 575) begin
					state<=2;
					out<=138;
				end
				if(in == 576) begin
					state<=2;
					out<=139;
				end
				if(in == 577) begin
					state<=2;
					out<=140;
				end
				if(in == 578) begin
					state<=2;
					out<=141;
				end
				if(in == 579) begin
					state<=2;
					out<=142;
				end
				if(in == 580) begin
					state<=2;
					out<=143;
				end
				if(in == 581) begin
					state<=3;
					out<=144;
				end
				if(in == 582) begin
					state<=11;
					out<=145;
				end
				if(in == 583) begin
					state<=3;
					out<=146;
				end
				if(in == 584) begin
					state<=12;
					out<=147;
				end
				if(in == 585) begin
					state<=3;
					out<=148;
				end
				if(in == 586) begin
					state<=12;
					out<=149;
				end
				if(in == 587) begin
					state<=12;
					out<=150;
				end
				if(in == 588) begin
					state<=12;
					out<=151;
				end
				if(in == 589) begin
					state<=12;
					out<=152;
				end
				if(in == 590) begin
					state<=12;
					out<=153;
				end
				if(in == 591) begin
					state<=12;
					out<=154;
				end
				if(in == 592) begin
					state<=12;
					out<=155;
				end
				if(in == 593) begin
					state<=12;
					out<=156;
				end
				if(in == 594) begin
					state<=12;
					out<=157;
				end
				if(in == 595) begin
					state<=12;
					out<=158;
				end
				if(in == 596) begin
					state<=12;
					out<=159;
				end
				if(in == 597) begin
					state<=12;
					out<=160;
				end
				if(in == 598) begin
					state<=12;
					out<=161;
				end
				if(in == 599) begin
					state<=12;
					out<=162;
				end
				if(in == 600) begin
					state<=12;
					out<=163;
				end
				if(in == 601) begin
					state<=12;
					out<=164;
				end
				if(in == 602) begin
					state<=12;
					out<=165;
				end
				if(in == 603) begin
					state<=12;
					out<=166;
				end
				if(in == 604) begin
					state<=12;
					out<=167;
				end
				if(in == 605) begin
					state<=12;
					out<=168;
				end
				if(in == 606) begin
					state<=12;
					out<=169;
				end
				if(in == 607) begin
					state<=12;
					out<=170;
				end
				if(in == 608) begin
					state<=12;
					out<=171;
				end
				if(in == 609) begin
					state<=12;
					out<=172;
				end
				if(in == 610) begin
					state<=12;
					out<=173;
				end
				if(in == 611) begin
					state<=12;
					out<=174;
				end
				if(in == 612) begin
					state<=12;
					out<=175;
				end
				if(in == 613) begin
					state<=12;
					out<=176;
				end
				if(in == 614) begin
					state<=12;
					out<=177;
				end
				if(in == 615) begin
					state<=12;
					out<=178;
				end
				if(in == 616) begin
					state<=12;
					out<=179;
				end
				if(in == 617) begin
					state<=12;
					out<=180;
				end
				if(in == 618) begin
					state<=12;
					out<=181;
				end
				if(in == 619) begin
					state<=12;
					out<=182;
				end
				if(in == 620) begin
					state<=12;
					out<=183;
				end
				if(in == 621) begin
					state<=12;
					out<=184;
				end
				if(in == 622) begin
					state<=12;
					out<=185;
				end
				if(in == 623) begin
					state<=12;
					out<=186;
				end
				if(in == 624) begin
					state<=12;
					out<=187;
				end
				if(in == 625) begin
					state<=12;
					out<=188;
				end
				if(in == 626) begin
					state<=12;
					out<=189;
				end
				if(in == 627) begin
					state<=12;
					out<=190;
				end
				if(in == 628) begin
					state<=12;
					out<=191;
				end
				if(in == 629) begin
					state<=12;
					out<=192;
				end
				if(in == 630) begin
					state<=12;
					out<=193;
				end
				if(in == 631) begin
					state<=12;
					out<=194;
				end
				if(in == 632) begin
					state<=12;
					out<=195;
				end
				if(in == 633) begin
					state<=3;
					out<=196;
				end
				if(in == 634) begin
					state<=11;
					out<=197;
				end
				if(in == 635) begin
					state<=3;
					out<=198;
				end
				if(in == 636) begin
					state<=12;
					out<=199;
				end
				if(in == 637) begin
					state<=3;
					out<=200;
				end
				if(in == 638) begin
					state<=12;
					out<=201;
				end
				if(in == 639) begin
					state<=12;
					out<=202;
				end
				if(in == 640) begin
					state<=12;
					out<=203;
				end
				if(in == 641) begin
					state<=12;
					out<=204;
				end
				if(in == 642) begin
					state<=12;
					out<=205;
				end
				if(in == 643) begin
					state<=12;
					out<=206;
				end
				if(in == 644) begin
					state<=12;
					out<=207;
				end
				if(in == 645) begin
					state<=12;
					out<=208;
				end
				if(in == 646) begin
					state<=12;
					out<=209;
				end
				if(in == 647) begin
					state<=12;
					out<=210;
				end
				if(in == 648) begin
					state<=12;
					out<=211;
				end
				if(in == 649) begin
					state<=12;
					out<=212;
				end
				if(in == 650) begin
					state<=12;
					out<=213;
				end
				if(in == 651) begin
					state<=12;
					out<=214;
				end
				if(in == 652) begin
					state<=12;
					out<=215;
				end
				if(in == 653) begin
					state<=12;
					out<=216;
				end
				if(in == 654) begin
					state<=12;
					out<=217;
				end
				if(in == 655) begin
					state<=12;
					out<=218;
				end
				if(in == 656) begin
					state<=12;
					out<=219;
				end
				if(in == 657) begin
					state<=12;
					out<=220;
				end
				if(in == 658) begin
					state<=12;
					out<=221;
				end
				if(in == 659) begin
					state<=12;
					out<=222;
				end
				if(in == 660) begin
					state<=12;
					out<=223;
				end
				if(in == 661) begin
					state<=12;
					out<=224;
				end
				if(in == 662) begin
					state<=12;
					out<=225;
				end
				if(in == 663) begin
					state<=12;
					out<=226;
				end
				if(in == 664) begin
					state<=12;
					out<=227;
				end
				if(in == 665) begin
					state<=12;
					out<=228;
				end
				if(in == 666) begin
					state<=12;
					out<=229;
				end
				if(in == 667) begin
					state<=12;
					out<=230;
				end
				if(in == 668) begin
					state<=12;
					out<=231;
				end
				if(in == 669) begin
					state<=12;
					out<=232;
				end
				if(in == 670) begin
					state<=12;
					out<=233;
				end
				if(in == 671) begin
					state<=12;
					out<=234;
				end
				if(in == 672) begin
					state<=12;
					out<=235;
				end
				if(in == 673) begin
					state<=12;
					out<=236;
				end
				if(in == 674) begin
					state<=12;
					out<=237;
				end
				if(in == 675) begin
					state<=12;
					out<=238;
				end
				if(in == 676) begin
					state<=12;
					out<=239;
				end
				if(in == 677) begin
					state<=12;
					out<=240;
				end
				if(in == 678) begin
					state<=12;
					out<=241;
				end
				if(in == 679) begin
					state<=12;
					out<=242;
				end
				if(in == 680) begin
					state<=12;
					out<=243;
				end
				if(in == 681) begin
					state<=12;
					out<=244;
				end
				if(in == 682) begin
					state<=12;
					out<=245;
				end
				if(in == 683) begin
					state<=12;
					out<=246;
				end
				if(in == 684) begin
					state<=12;
					out<=247;
				end
				if(in == 685) begin
					state<=2;
					out<=248;
				end
				if(in == 686) begin
					state<=2;
					out<=249;
				end
				if(in == 687) begin
					state<=2;
					out<=250;
				end
				if(in == 688) begin
					state<=2;
					out<=251;
				end
				if(in == 689) begin
					state<=2;
					out<=252;
				end
				if(in == 690) begin
					state<=2;
					out<=253;
				end
				if(in == 691) begin
					state<=2;
					out<=254;
				end
				if(in == 692) begin
					state<=2;
					out<=255;
				end
				if(in == 693) begin
					state<=2;
					out<=0;
				end
				if(in == 694) begin
					state<=2;
					out<=1;
				end
				if(in == 695) begin
					state<=2;
					out<=2;
				end
				if(in == 696) begin
					state<=2;
					out<=3;
				end
				if(in == 697) begin
					state<=3;
					out<=4;
				end
				if(in == 698) begin
					state<=11;
					out<=5;
				end
				if(in == 699) begin
					state<=3;
					out<=6;
				end
				if(in == 700) begin
					state<=12;
					out<=7;
				end
				if(in == 701) begin
					state<=3;
					out<=8;
				end
				if(in == 702) begin
					state<=12;
					out<=9;
				end
				if(in == 703) begin
					state<=12;
					out<=10;
				end
				if(in == 704) begin
					state<=12;
					out<=11;
				end
				if(in == 705) begin
					state<=12;
					out<=12;
				end
				if(in == 706) begin
					state<=12;
					out<=13;
				end
				if(in == 707) begin
					state<=12;
					out<=14;
				end
				if(in == 708) begin
					state<=12;
					out<=15;
				end
				if(in == 709) begin
					state<=12;
					out<=16;
				end
				if(in == 710) begin
					state<=12;
					out<=17;
				end
				if(in == 711) begin
					state<=12;
					out<=18;
				end
				if(in == 712) begin
					state<=12;
					out<=19;
				end
				if(in == 713) begin
					state<=12;
					out<=20;
				end
				if(in == 714) begin
					state<=12;
					out<=21;
				end
				if(in == 715) begin
					state<=12;
					out<=22;
				end
				if(in == 716) begin
					state<=12;
					out<=23;
				end
				if(in == 717) begin
					state<=12;
					out<=24;
				end
				if(in == 718) begin
					state<=12;
					out<=25;
				end
				if(in == 719) begin
					state<=12;
					out<=26;
				end
				if(in == 720) begin
					state<=12;
					out<=27;
				end
				if(in == 721) begin
					state<=12;
					out<=28;
				end
				if(in == 722) begin
					state<=12;
					out<=29;
				end
				if(in == 723) begin
					state<=12;
					out<=30;
				end
				if(in == 724) begin
					state<=12;
					out<=31;
				end
				if(in == 725) begin
					state<=12;
					out<=32;
				end
				if(in == 726) begin
					state<=12;
					out<=33;
				end
				if(in == 727) begin
					state<=12;
					out<=34;
				end
				if(in == 728) begin
					state<=12;
					out<=35;
				end
				if(in == 729) begin
					state<=12;
					out<=36;
				end
				if(in == 730) begin
					state<=12;
					out<=37;
				end
				if(in == 731) begin
					state<=12;
					out<=38;
				end
				if(in == 732) begin
					state<=12;
					out<=39;
				end
				if(in == 733) begin
					state<=12;
					out<=40;
				end
				if(in == 734) begin
					state<=12;
					out<=41;
				end
				if(in == 735) begin
					state<=12;
					out<=42;
				end
				if(in == 736) begin
					state<=12;
					out<=43;
				end
				if(in == 737) begin
					state<=12;
					out<=44;
				end
				if(in == 738) begin
					state<=12;
					out<=45;
				end
				if(in == 739) begin
					state<=12;
					out<=46;
				end
				if(in == 740) begin
					state<=12;
					out<=47;
				end
				if(in == 741) begin
					state<=12;
					out<=48;
				end
				if(in == 742) begin
					state<=12;
					out<=49;
				end
				if(in == 743) begin
					state<=12;
					out<=50;
				end
				if(in == 744) begin
					state<=12;
					out<=51;
				end
				if(in == 745) begin
					state<=12;
					out<=52;
				end
				if(in == 746) begin
					state<=12;
					out<=53;
				end
				if(in == 747) begin
					state<=12;
					out<=54;
				end
				if(in == 748) begin
					state<=12;
					out<=55;
				end
				if(in == 749) begin
					state<=3;
					out<=56;
				end
				if(in == 750) begin
					state<=11;
					out<=57;
				end
				if(in == 751) begin
					state<=3;
					out<=58;
				end
				if(in == 752) begin
					state<=12;
					out<=59;
				end
				if(in == 753) begin
					state<=3;
					out<=60;
				end
				if(in == 754) begin
					state<=12;
					out<=61;
				end
				if(in == 755) begin
					state<=12;
					out<=62;
				end
				if(in == 756) begin
					state<=12;
					out<=63;
				end
				if(in == 757) begin
					state<=12;
					out<=64;
				end
				if(in == 758) begin
					state<=12;
					out<=65;
				end
				if(in == 759) begin
					state<=12;
					out<=66;
				end
				if(in == 760) begin
					state<=12;
					out<=67;
				end
				if(in == 761) begin
					state<=12;
					out<=68;
				end
				if(in == 762) begin
					state<=12;
					out<=69;
				end
				if(in == 763) begin
					state<=12;
					out<=70;
				end
				if(in == 764) begin
					state<=12;
					out<=71;
				end
				if(in == 765) begin
					state<=12;
					out<=72;
				end
				if(in == 766) begin
					state<=12;
					out<=73;
				end
				if(in == 767) begin
					state<=12;
					out<=74;
				end
				if(in == 768) begin
					state<=12;
					out<=75;
				end
				if(in == 769) begin
					state<=12;
					out<=76;
				end
				if(in == 770) begin
					state<=12;
					out<=77;
				end
				if(in == 771) begin
					state<=12;
					out<=78;
				end
				if(in == 772) begin
					state<=12;
					out<=79;
				end
				if(in == 773) begin
					state<=12;
					out<=80;
				end
				if(in == 774) begin
					state<=12;
					out<=81;
				end
				if(in == 775) begin
					state<=12;
					out<=82;
				end
				if(in == 776) begin
					state<=12;
					out<=83;
				end
				if(in == 777) begin
					state<=12;
					out<=84;
				end
				if(in == 778) begin
					state<=12;
					out<=85;
				end
				if(in == 779) begin
					state<=12;
					out<=86;
				end
				if(in == 780) begin
					state<=12;
					out<=87;
				end
				if(in == 781) begin
					state<=12;
					out<=88;
				end
				if(in == 782) begin
					state<=12;
					out<=89;
				end
				if(in == 783) begin
					state<=12;
					out<=90;
				end
				if(in == 784) begin
					state<=12;
					out<=91;
				end
				if(in == 785) begin
					state<=12;
					out<=92;
				end
				if(in == 786) begin
					state<=12;
					out<=93;
				end
				if(in == 787) begin
					state<=12;
					out<=94;
				end
				if(in == 788) begin
					state<=12;
					out<=95;
				end
				if(in == 789) begin
					state<=12;
					out<=96;
				end
				if(in == 790) begin
					state<=12;
					out<=97;
				end
				if(in == 791) begin
					state<=12;
					out<=98;
				end
				if(in == 792) begin
					state<=12;
					out<=99;
				end
				if(in == 793) begin
					state<=12;
					out<=100;
				end
				if(in == 794) begin
					state<=12;
					out<=101;
				end
				if(in == 795) begin
					state<=12;
					out<=102;
				end
				if(in == 796) begin
					state<=12;
					out<=103;
				end
				if(in == 797) begin
					state<=12;
					out<=104;
				end
				if(in == 798) begin
					state<=12;
					out<=105;
				end
				if(in == 799) begin
					state<=12;
					out<=106;
				end
				if(in == 800) begin
					state<=12;
					out<=107;
				end
				if(in == 801) begin
					state<=2;
					out<=108;
				end
				if(in == 802) begin
					state<=2;
					out<=109;
				end
				if(in == 803) begin
					state<=2;
					out<=110;
				end
				if(in == 804) begin
					state<=2;
					out<=111;
				end
				if(in == 805) begin
					state<=2;
					out<=112;
				end
				if(in == 806) begin
					state<=2;
					out<=113;
				end
				if(in == 807) begin
					state<=2;
					out<=114;
				end
				if(in == 808) begin
					state<=2;
					out<=115;
				end
				if(in == 809) begin
					state<=2;
					out<=116;
				end
				if(in == 810) begin
					state<=2;
					out<=117;
				end
				if(in == 811) begin
					state<=2;
					out<=118;
				end
				if(in == 812) begin
					state<=2;
					out<=119;
				end
				if(in == 813) begin
					state<=3;
					out<=120;
				end
				if(in == 814) begin
					state<=11;
					out<=121;
				end
				if(in == 815) begin
					state<=3;
					out<=122;
				end
				if(in == 816) begin
					state<=12;
					out<=123;
				end
				if(in == 817) begin
					state<=3;
					out<=124;
				end
				if(in == 818) begin
					state<=12;
					out<=125;
				end
				if(in == 819) begin
					state<=12;
					out<=126;
				end
				if(in == 820) begin
					state<=12;
					out<=127;
				end
				if(in == 821) begin
					state<=12;
					out<=128;
				end
				if(in == 822) begin
					state<=12;
					out<=129;
				end
				if(in == 823) begin
					state<=12;
					out<=130;
				end
				if(in == 824) begin
					state<=12;
					out<=131;
				end
				if(in == 825) begin
					state<=12;
					out<=132;
				end
				if(in == 826) begin
					state<=12;
					out<=133;
				end
				if(in == 827) begin
					state<=12;
					out<=134;
				end
				if(in == 828) begin
					state<=12;
					out<=135;
				end
				if(in == 829) begin
					state<=12;
					out<=136;
				end
				if(in == 830) begin
					state<=12;
					out<=137;
				end
				if(in == 831) begin
					state<=12;
					out<=138;
				end
				if(in == 832) begin
					state<=12;
					out<=139;
				end
				if(in == 833) begin
					state<=12;
					out<=140;
				end
				if(in == 834) begin
					state<=12;
					out<=141;
				end
				if(in == 835) begin
					state<=12;
					out<=142;
				end
				if(in == 836) begin
					state<=12;
					out<=143;
				end
				if(in == 837) begin
					state<=12;
					out<=144;
				end
				if(in == 838) begin
					state<=12;
					out<=145;
				end
				if(in == 839) begin
					state<=12;
					out<=146;
				end
				if(in == 840) begin
					state<=12;
					out<=147;
				end
				if(in == 841) begin
					state<=12;
					out<=148;
				end
				if(in == 842) begin
					state<=12;
					out<=149;
				end
				if(in == 843) begin
					state<=12;
					out<=150;
				end
				if(in == 844) begin
					state<=12;
					out<=151;
				end
				if(in == 845) begin
					state<=12;
					out<=152;
				end
				if(in == 846) begin
					state<=12;
					out<=153;
				end
				if(in == 847) begin
					state<=12;
					out<=154;
				end
				if(in == 848) begin
					state<=12;
					out<=155;
				end
				if(in == 849) begin
					state<=12;
					out<=156;
				end
				if(in == 850) begin
					state<=12;
					out<=157;
				end
				if(in == 851) begin
					state<=12;
					out<=158;
				end
				if(in == 852) begin
					state<=12;
					out<=159;
				end
				if(in == 853) begin
					state<=12;
					out<=160;
				end
				if(in == 854) begin
					state<=12;
					out<=161;
				end
				if(in == 855) begin
					state<=12;
					out<=162;
				end
				if(in == 856) begin
					state<=12;
					out<=163;
				end
				if(in == 857) begin
					state<=12;
					out<=164;
				end
				if(in == 858) begin
					state<=12;
					out<=165;
				end
				if(in == 859) begin
					state<=12;
					out<=166;
				end
				if(in == 860) begin
					state<=12;
					out<=167;
				end
				if(in == 861) begin
					state<=12;
					out<=168;
				end
				if(in == 862) begin
					state<=12;
					out<=169;
				end
				if(in == 863) begin
					state<=12;
					out<=170;
				end
				if(in == 864) begin
					state<=12;
					out<=171;
				end
				if(in == 865) begin
					state<=3;
					out<=172;
				end
				if(in == 866) begin
					state<=11;
					out<=173;
				end
				if(in == 867) begin
					state<=3;
					out<=174;
				end
				if(in == 868) begin
					state<=12;
					out<=175;
				end
				if(in == 869) begin
					state<=3;
					out<=176;
				end
				if(in == 870) begin
					state<=12;
					out<=177;
				end
				if(in == 871) begin
					state<=12;
					out<=178;
				end
				if(in == 872) begin
					state<=12;
					out<=179;
				end
				if(in == 873) begin
					state<=12;
					out<=180;
				end
				if(in == 874) begin
					state<=12;
					out<=181;
				end
				if(in == 875) begin
					state<=12;
					out<=182;
				end
				if(in == 876) begin
					state<=12;
					out<=183;
				end
				if(in == 877) begin
					state<=12;
					out<=184;
				end
				if(in == 878) begin
					state<=12;
					out<=185;
				end
				if(in == 879) begin
					state<=12;
					out<=186;
				end
				if(in == 880) begin
					state<=12;
					out<=187;
				end
				if(in == 881) begin
					state<=12;
					out<=188;
				end
				if(in == 882) begin
					state<=12;
					out<=189;
				end
				if(in == 883) begin
					state<=12;
					out<=190;
				end
				if(in == 884) begin
					state<=12;
					out<=191;
				end
				if(in == 885) begin
					state<=12;
					out<=192;
				end
				if(in == 886) begin
					state<=12;
					out<=193;
				end
				if(in == 887) begin
					state<=12;
					out<=194;
				end
				if(in == 888) begin
					state<=12;
					out<=195;
				end
				if(in == 889) begin
					state<=12;
					out<=196;
				end
				if(in == 890) begin
					state<=12;
					out<=197;
				end
				if(in == 891) begin
					state<=12;
					out<=198;
				end
				if(in == 892) begin
					state<=12;
					out<=199;
				end
				if(in == 893) begin
					state<=12;
					out<=200;
				end
				if(in == 894) begin
					state<=12;
					out<=201;
				end
				if(in == 895) begin
					state<=12;
					out<=202;
				end
				if(in == 896) begin
					state<=12;
					out<=203;
				end
				if(in == 897) begin
					state<=12;
					out<=204;
				end
				if(in == 898) begin
					state<=12;
					out<=205;
				end
				if(in == 899) begin
					state<=12;
					out<=206;
				end
				if(in == 900) begin
					state<=12;
					out<=207;
				end
				if(in == 901) begin
					state<=12;
					out<=208;
				end
				if(in == 902) begin
					state<=12;
					out<=209;
				end
				if(in == 903) begin
					state<=12;
					out<=210;
				end
				if(in == 904) begin
					state<=12;
					out<=211;
				end
				if(in == 905) begin
					state<=12;
					out<=212;
				end
				if(in == 906) begin
					state<=12;
					out<=213;
				end
				if(in == 907) begin
					state<=12;
					out<=214;
				end
				if(in == 908) begin
					state<=12;
					out<=215;
				end
				if(in == 909) begin
					state<=12;
					out<=216;
				end
				if(in == 910) begin
					state<=12;
					out<=217;
				end
				if(in == 911) begin
					state<=12;
					out<=218;
				end
				if(in == 912) begin
					state<=12;
					out<=219;
				end
				if(in == 913) begin
					state<=12;
					out<=220;
				end
				if(in == 914) begin
					state<=12;
					out<=221;
				end
				if(in == 915) begin
					state<=12;
					out<=222;
				end
				if(in == 916) begin
					state<=12;
					out<=223;
				end
				if(in == 917) begin
					state<=2;
					out<=224;
				end
				if(in == 918) begin
					state<=2;
					out<=225;
				end
				if(in == 919) begin
					state<=2;
					out<=226;
				end
				if(in == 920) begin
					state<=2;
					out<=227;
				end
				if(in == 921) begin
					state<=2;
					out<=228;
				end
				if(in == 922) begin
					state<=2;
					out<=229;
				end
				if(in == 923) begin
					state<=2;
					out<=230;
				end
				if(in == 924) begin
					state<=2;
					out<=231;
				end
				if(in == 925) begin
					state<=2;
					out<=232;
				end
				if(in == 926) begin
					state<=2;
					out<=233;
				end
				if(in == 927) begin
					state<=2;
					out<=234;
				end
				if(in == 928) begin
					state<=2;
					out<=235;
				end
			end
			12: begin
				if(in == 0) begin
					state<=13;
					out<=236;
				end
				if(in == 1) begin
					state<=1;
					out<=237;
				end
				if(in == 2) begin
					state<=12;
					out<=238;
				end
				if(in == 3) begin
					state<=13;
					out<=239;
				end
				if(in == 4) begin
					state<=12;
					out<=240;
				end
				if(in == 5) begin
					state<=13;
					out<=241;
				end
				if(in == 6) begin
					state<=12;
					out<=242;
				end
				if(in == 7) begin
					state<=12;
					out<=243;
				end
				if(in == 8) begin
					state<=12;
					out<=244;
				end
				if(in == 9) begin
					state<=12;
					out<=245;
				end
				if(in == 10) begin
					state<=12;
					out<=246;
				end
				if(in == 11) begin
					state<=12;
					out<=247;
				end
				if(in == 12) begin
					state<=12;
					out<=248;
				end
				if(in == 13) begin
					state<=12;
					out<=249;
				end
				if(in == 14) begin
					state<=12;
					out<=250;
				end
				if(in == 15) begin
					state<=12;
					out<=251;
				end
				if(in == 16) begin
					state<=12;
					out<=252;
				end
				if(in == 17) begin
					state<=12;
					out<=253;
				end
				if(in == 18) begin
					state<=12;
					out<=254;
				end
				if(in == 19) begin
					state<=12;
					out<=255;
				end
				if(in == 20) begin
					state<=12;
					out<=0;
				end
				if(in == 21) begin
					state<=12;
					out<=1;
				end
				if(in == 22) begin
					state<=12;
					out<=2;
				end
				if(in == 23) begin
					state<=12;
					out<=3;
				end
				if(in == 24) begin
					state<=12;
					out<=4;
				end
				if(in == 25) begin
					state<=12;
					out<=5;
				end
				if(in == 26) begin
					state<=12;
					out<=6;
				end
				if(in == 27) begin
					state<=12;
					out<=7;
				end
				if(in == 28) begin
					state<=12;
					out<=8;
				end
				if(in == 29) begin
					state<=12;
					out<=9;
				end
				if(in == 30) begin
					state<=12;
					out<=10;
				end
				if(in == 31) begin
					state<=12;
					out<=11;
				end
				if(in == 32) begin
					state<=12;
					out<=12;
				end
				if(in == 33) begin
					state<=12;
					out<=13;
				end
				if(in == 34) begin
					state<=12;
					out<=14;
				end
				if(in == 35) begin
					state<=12;
					out<=15;
				end
				if(in == 36) begin
					state<=12;
					out<=16;
				end
				if(in == 37) begin
					state<=12;
					out<=17;
				end
				if(in == 38) begin
					state<=12;
					out<=18;
				end
				if(in == 39) begin
					state<=12;
					out<=19;
				end
				if(in == 40) begin
					state<=12;
					out<=20;
				end
				if(in == 41) begin
					state<=12;
					out<=21;
				end
				if(in == 42) begin
					state<=12;
					out<=22;
				end
				if(in == 43) begin
					state<=12;
					out<=23;
				end
				if(in == 44) begin
					state<=12;
					out<=24;
				end
				if(in == 45) begin
					state<=12;
					out<=25;
				end
				if(in == 46) begin
					state<=12;
					out<=26;
				end
				if(in == 47) begin
					state<=12;
					out<=27;
				end
				if(in == 48) begin
					state<=12;
					out<=28;
				end
				if(in == 49) begin
					state<=12;
					out<=29;
				end
				if(in == 50) begin
					state<=12;
					out<=30;
				end
				if(in == 51) begin
					state<=12;
					out<=31;
				end
				if(in == 52) begin
					state<=12;
					out<=32;
				end
				if(in == 53) begin
					state<=13;
					out<=33;
				end
				if(in == 54) begin
					state<=12;
					out<=34;
				end
				if(in == 55) begin
					state<=13;
					out<=35;
				end
				if(in == 56) begin
					state<=12;
					out<=36;
				end
				if(in == 57) begin
					state<=13;
					out<=37;
				end
				if(in == 58) begin
					state<=12;
					out<=38;
				end
				if(in == 59) begin
					state<=12;
					out<=39;
				end
				if(in == 60) begin
					state<=12;
					out<=40;
				end
				if(in == 61) begin
					state<=12;
					out<=41;
				end
				if(in == 62) begin
					state<=12;
					out<=42;
				end
				if(in == 63) begin
					state<=12;
					out<=43;
				end
				if(in == 64) begin
					state<=12;
					out<=44;
				end
				if(in == 65) begin
					state<=12;
					out<=45;
				end
				if(in == 66) begin
					state<=12;
					out<=46;
				end
				if(in == 67) begin
					state<=12;
					out<=47;
				end
				if(in == 68) begin
					state<=12;
					out<=48;
				end
				if(in == 69) begin
					state<=12;
					out<=49;
				end
				if(in == 70) begin
					state<=12;
					out<=50;
				end
				if(in == 71) begin
					state<=12;
					out<=51;
				end
				if(in == 72) begin
					state<=12;
					out<=52;
				end
				if(in == 73) begin
					state<=12;
					out<=53;
				end
				if(in == 74) begin
					state<=12;
					out<=54;
				end
				if(in == 75) begin
					state<=12;
					out<=55;
				end
				if(in == 76) begin
					state<=12;
					out<=56;
				end
				if(in == 77) begin
					state<=12;
					out<=57;
				end
				if(in == 78) begin
					state<=12;
					out<=58;
				end
				if(in == 79) begin
					state<=12;
					out<=59;
				end
				if(in == 80) begin
					state<=12;
					out<=60;
				end
				if(in == 81) begin
					state<=12;
					out<=61;
				end
				if(in == 82) begin
					state<=12;
					out<=62;
				end
				if(in == 83) begin
					state<=12;
					out<=63;
				end
				if(in == 84) begin
					state<=12;
					out<=64;
				end
				if(in == 85) begin
					state<=12;
					out<=65;
				end
				if(in == 86) begin
					state<=12;
					out<=66;
				end
				if(in == 87) begin
					state<=12;
					out<=67;
				end
				if(in == 88) begin
					state<=12;
					out<=68;
				end
				if(in == 89) begin
					state<=12;
					out<=69;
				end
				if(in == 90) begin
					state<=12;
					out<=70;
				end
				if(in == 91) begin
					state<=12;
					out<=71;
				end
				if(in == 92) begin
					state<=12;
					out<=72;
				end
				if(in == 93) begin
					state<=12;
					out<=73;
				end
				if(in == 94) begin
					state<=12;
					out<=74;
				end
				if(in == 95) begin
					state<=12;
					out<=75;
				end
				if(in == 96) begin
					state<=12;
					out<=76;
				end
				if(in == 97) begin
					state<=12;
					out<=77;
				end
				if(in == 98) begin
					state<=12;
					out<=78;
				end
				if(in == 99) begin
					state<=12;
					out<=79;
				end
				if(in == 100) begin
					state<=12;
					out<=80;
				end
				if(in == 101) begin
					state<=12;
					out<=81;
				end
				if(in == 102) begin
					state<=12;
					out<=82;
				end
				if(in == 103) begin
					state<=12;
					out<=83;
				end
				if(in == 104) begin
					state<=12;
					out<=84;
				end
				if(in == 105) begin
					state<=2;
					out<=85;
				end
				if(in == 106) begin
					state<=2;
					out<=86;
				end
				if(in == 107) begin
					state<=2;
					out<=87;
				end
				if(in == 108) begin
					state<=2;
					out<=88;
				end
				if(in == 109) begin
					state<=2;
					out<=89;
				end
				if(in == 110) begin
					state<=2;
					out<=90;
				end
				if(in == 111) begin
					state<=2;
					out<=91;
				end
				if(in == 112) begin
					state<=2;
					out<=92;
				end
				if(in == 113) begin
					state<=2;
					out<=93;
				end
				if(in == 114) begin
					state<=2;
					out<=94;
				end
				if(in == 115) begin
					state<=2;
					out<=95;
				end
				if(in == 116) begin
					state<=2;
					out<=96;
				end
				if(in == 117) begin
					state<=13;
					out<=97;
				end
				if(in == 118) begin
					state<=12;
					out<=98;
				end
				if(in == 119) begin
					state<=13;
					out<=99;
				end
				if(in == 120) begin
					state<=12;
					out<=100;
				end
				if(in == 121) begin
					state<=13;
					out<=101;
				end
				if(in == 122) begin
					state<=12;
					out<=102;
				end
				if(in == 123) begin
					state<=12;
					out<=103;
				end
				if(in == 124) begin
					state<=12;
					out<=104;
				end
				if(in == 125) begin
					state<=12;
					out<=105;
				end
				if(in == 126) begin
					state<=12;
					out<=106;
				end
				if(in == 127) begin
					state<=12;
					out<=107;
				end
				if(in == 128) begin
					state<=12;
					out<=108;
				end
				if(in == 129) begin
					state<=12;
					out<=109;
				end
				if(in == 130) begin
					state<=12;
					out<=110;
				end
				if(in == 131) begin
					state<=12;
					out<=111;
				end
				if(in == 132) begin
					state<=12;
					out<=112;
				end
				if(in == 133) begin
					state<=12;
					out<=113;
				end
				if(in == 134) begin
					state<=12;
					out<=114;
				end
				if(in == 135) begin
					state<=12;
					out<=115;
				end
				if(in == 136) begin
					state<=12;
					out<=116;
				end
				if(in == 137) begin
					state<=12;
					out<=117;
				end
				if(in == 138) begin
					state<=12;
					out<=118;
				end
				if(in == 139) begin
					state<=12;
					out<=119;
				end
				if(in == 140) begin
					state<=12;
					out<=120;
				end
				if(in == 141) begin
					state<=12;
					out<=121;
				end
				if(in == 142) begin
					state<=12;
					out<=122;
				end
				if(in == 143) begin
					state<=12;
					out<=123;
				end
				if(in == 144) begin
					state<=12;
					out<=124;
				end
				if(in == 145) begin
					state<=12;
					out<=125;
				end
				if(in == 146) begin
					state<=12;
					out<=126;
				end
				if(in == 147) begin
					state<=12;
					out<=127;
				end
				if(in == 148) begin
					state<=12;
					out<=128;
				end
				if(in == 149) begin
					state<=12;
					out<=129;
				end
				if(in == 150) begin
					state<=12;
					out<=130;
				end
				if(in == 151) begin
					state<=12;
					out<=131;
				end
				if(in == 152) begin
					state<=12;
					out<=132;
				end
				if(in == 153) begin
					state<=12;
					out<=133;
				end
				if(in == 154) begin
					state<=12;
					out<=134;
				end
				if(in == 155) begin
					state<=12;
					out<=135;
				end
				if(in == 156) begin
					state<=12;
					out<=136;
				end
				if(in == 157) begin
					state<=12;
					out<=137;
				end
				if(in == 158) begin
					state<=12;
					out<=138;
				end
				if(in == 159) begin
					state<=12;
					out<=139;
				end
				if(in == 160) begin
					state<=12;
					out<=140;
				end
				if(in == 161) begin
					state<=12;
					out<=141;
				end
				if(in == 162) begin
					state<=12;
					out<=142;
				end
				if(in == 163) begin
					state<=12;
					out<=143;
				end
				if(in == 164) begin
					state<=12;
					out<=144;
				end
				if(in == 165) begin
					state<=12;
					out<=145;
				end
				if(in == 166) begin
					state<=12;
					out<=146;
				end
				if(in == 167) begin
					state<=12;
					out<=147;
				end
				if(in == 168) begin
					state<=12;
					out<=148;
				end
				if(in == 169) begin
					state<=13;
					out<=149;
				end
				if(in == 170) begin
					state<=12;
					out<=150;
				end
				if(in == 171) begin
					state<=13;
					out<=151;
				end
				if(in == 172) begin
					state<=12;
					out<=152;
				end
				if(in == 173) begin
					state<=13;
					out<=153;
				end
				if(in == 174) begin
					state<=12;
					out<=154;
				end
				if(in == 175) begin
					state<=12;
					out<=155;
				end
				if(in == 176) begin
					state<=12;
					out<=156;
				end
				if(in == 177) begin
					state<=12;
					out<=157;
				end
				if(in == 178) begin
					state<=12;
					out<=158;
				end
				if(in == 179) begin
					state<=12;
					out<=159;
				end
				if(in == 180) begin
					state<=12;
					out<=160;
				end
				if(in == 181) begin
					state<=12;
					out<=161;
				end
				if(in == 182) begin
					state<=12;
					out<=162;
				end
				if(in == 183) begin
					state<=12;
					out<=163;
				end
				if(in == 184) begin
					state<=12;
					out<=164;
				end
				if(in == 185) begin
					state<=12;
					out<=165;
				end
				if(in == 186) begin
					state<=12;
					out<=166;
				end
				if(in == 187) begin
					state<=12;
					out<=167;
				end
				if(in == 188) begin
					state<=12;
					out<=168;
				end
				if(in == 189) begin
					state<=12;
					out<=169;
				end
				if(in == 190) begin
					state<=12;
					out<=170;
				end
				if(in == 191) begin
					state<=12;
					out<=171;
				end
				if(in == 192) begin
					state<=12;
					out<=172;
				end
				if(in == 193) begin
					state<=12;
					out<=173;
				end
				if(in == 194) begin
					state<=12;
					out<=174;
				end
				if(in == 195) begin
					state<=12;
					out<=175;
				end
				if(in == 196) begin
					state<=12;
					out<=176;
				end
				if(in == 197) begin
					state<=12;
					out<=177;
				end
				if(in == 198) begin
					state<=12;
					out<=178;
				end
				if(in == 199) begin
					state<=12;
					out<=179;
				end
				if(in == 200) begin
					state<=12;
					out<=180;
				end
				if(in == 201) begin
					state<=12;
					out<=181;
				end
				if(in == 202) begin
					state<=12;
					out<=182;
				end
				if(in == 203) begin
					state<=12;
					out<=183;
				end
				if(in == 204) begin
					state<=12;
					out<=184;
				end
				if(in == 205) begin
					state<=12;
					out<=185;
				end
				if(in == 206) begin
					state<=12;
					out<=186;
				end
				if(in == 207) begin
					state<=12;
					out<=187;
				end
				if(in == 208) begin
					state<=12;
					out<=188;
				end
				if(in == 209) begin
					state<=12;
					out<=189;
				end
				if(in == 210) begin
					state<=12;
					out<=190;
				end
				if(in == 211) begin
					state<=12;
					out<=191;
				end
				if(in == 212) begin
					state<=12;
					out<=192;
				end
				if(in == 213) begin
					state<=12;
					out<=193;
				end
				if(in == 214) begin
					state<=12;
					out<=194;
				end
				if(in == 215) begin
					state<=12;
					out<=195;
				end
				if(in == 216) begin
					state<=12;
					out<=196;
				end
				if(in == 217) begin
					state<=12;
					out<=197;
				end
				if(in == 218) begin
					state<=12;
					out<=198;
				end
				if(in == 219) begin
					state<=12;
					out<=199;
				end
				if(in == 220) begin
					state<=12;
					out<=200;
				end
				if(in == 221) begin
					state<=2;
					out<=201;
				end
				if(in == 222) begin
					state<=2;
					out<=202;
				end
				if(in == 223) begin
					state<=2;
					out<=203;
				end
				if(in == 224) begin
					state<=2;
					out<=204;
				end
				if(in == 225) begin
					state<=2;
					out<=205;
				end
				if(in == 226) begin
					state<=2;
					out<=206;
				end
				if(in == 227) begin
					state<=2;
					out<=207;
				end
				if(in == 228) begin
					state<=2;
					out<=208;
				end
				if(in == 229) begin
					state<=2;
					out<=209;
				end
				if(in == 230) begin
					state<=2;
					out<=210;
				end
				if(in == 231) begin
					state<=2;
					out<=211;
				end
				if(in == 232) begin
					state<=2;
					out<=212;
				end
				if(in == 233) begin
					state<=13;
					out<=213;
				end
				if(in == 234) begin
					state<=12;
					out<=214;
				end
				if(in == 235) begin
					state<=13;
					out<=215;
				end
				if(in == 236) begin
					state<=12;
					out<=216;
				end
				if(in == 237) begin
					state<=13;
					out<=217;
				end
				if(in == 238) begin
					state<=12;
					out<=218;
				end
				if(in == 239) begin
					state<=12;
					out<=219;
				end
				if(in == 240) begin
					state<=12;
					out<=220;
				end
				if(in == 241) begin
					state<=12;
					out<=221;
				end
				if(in == 242) begin
					state<=12;
					out<=222;
				end
				if(in == 243) begin
					state<=12;
					out<=223;
				end
				if(in == 244) begin
					state<=12;
					out<=224;
				end
				if(in == 245) begin
					state<=12;
					out<=225;
				end
				if(in == 246) begin
					state<=12;
					out<=226;
				end
				if(in == 247) begin
					state<=12;
					out<=227;
				end
				if(in == 248) begin
					state<=12;
					out<=228;
				end
				if(in == 249) begin
					state<=12;
					out<=229;
				end
				if(in == 250) begin
					state<=12;
					out<=230;
				end
				if(in == 251) begin
					state<=12;
					out<=231;
				end
				if(in == 252) begin
					state<=12;
					out<=232;
				end
				if(in == 253) begin
					state<=12;
					out<=233;
				end
				if(in == 254) begin
					state<=12;
					out<=234;
				end
				if(in == 255) begin
					state<=12;
					out<=235;
				end
				if(in == 256) begin
					state<=12;
					out<=236;
				end
				if(in == 257) begin
					state<=12;
					out<=237;
				end
				if(in == 258) begin
					state<=12;
					out<=238;
				end
				if(in == 259) begin
					state<=12;
					out<=239;
				end
				if(in == 260) begin
					state<=12;
					out<=240;
				end
				if(in == 261) begin
					state<=12;
					out<=241;
				end
				if(in == 262) begin
					state<=12;
					out<=242;
				end
				if(in == 263) begin
					state<=12;
					out<=243;
				end
				if(in == 264) begin
					state<=12;
					out<=244;
				end
				if(in == 265) begin
					state<=12;
					out<=245;
				end
				if(in == 266) begin
					state<=12;
					out<=246;
				end
				if(in == 267) begin
					state<=12;
					out<=247;
				end
				if(in == 268) begin
					state<=12;
					out<=248;
				end
				if(in == 269) begin
					state<=12;
					out<=249;
				end
				if(in == 270) begin
					state<=12;
					out<=250;
				end
				if(in == 271) begin
					state<=12;
					out<=251;
				end
				if(in == 272) begin
					state<=12;
					out<=252;
				end
				if(in == 273) begin
					state<=12;
					out<=253;
				end
				if(in == 274) begin
					state<=12;
					out<=254;
				end
				if(in == 275) begin
					state<=12;
					out<=255;
				end
				if(in == 276) begin
					state<=12;
					out<=0;
				end
				if(in == 277) begin
					state<=12;
					out<=1;
				end
				if(in == 278) begin
					state<=12;
					out<=2;
				end
				if(in == 279) begin
					state<=12;
					out<=3;
				end
				if(in == 280) begin
					state<=12;
					out<=4;
				end
				if(in == 281) begin
					state<=12;
					out<=5;
				end
				if(in == 282) begin
					state<=12;
					out<=6;
				end
				if(in == 283) begin
					state<=12;
					out<=7;
				end
				if(in == 284) begin
					state<=12;
					out<=8;
				end
				if(in == 285) begin
					state<=13;
					out<=9;
				end
				if(in == 286) begin
					state<=12;
					out<=10;
				end
				if(in == 287) begin
					state<=13;
					out<=11;
				end
				if(in == 288) begin
					state<=12;
					out<=12;
				end
				if(in == 289) begin
					state<=13;
					out<=13;
				end
				if(in == 290) begin
					state<=12;
					out<=14;
				end
				if(in == 291) begin
					state<=12;
					out<=15;
				end
				if(in == 292) begin
					state<=12;
					out<=16;
				end
				if(in == 293) begin
					state<=12;
					out<=17;
				end
				if(in == 294) begin
					state<=12;
					out<=18;
				end
				if(in == 295) begin
					state<=12;
					out<=19;
				end
				if(in == 296) begin
					state<=12;
					out<=20;
				end
				if(in == 297) begin
					state<=12;
					out<=21;
				end
				if(in == 298) begin
					state<=12;
					out<=22;
				end
				if(in == 299) begin
					state<=12;
					out<=23;
				end
				if(in == 300) begin
					state<=12;
					out<=24;
				end
				if(in == 301) begin
					state<=12;
					out<=25;
				end
				if(in == 302) begin
					state<=12;
					out<=26;
				end
				if(in == 303) begin
					state<=12;
					out<=27;
				end
				if(in == 304) begin
					state<=12;
					out<=28;
				end
				if(in == 305) begin
					state<=12;
					out<=29;
				end
				if(in == 306) begin
					state<=12;
					out<=30;
				end
				if(in == 307) begin
					state<=12;
					out<=31;
				end
				if(in == 308) begin
					state<=12;
					out<=32;
				end
				if(in == 309) begin
					state<=12;
					out<=33;
				end
				if(in == 310) begin
					state<=12;
					out<=34;
				end
				if(in == 311) begin
					state<=12;
					out<=35;
				end
				if(in == 312) begin
					state<=12;
					out<=36;
				end
				if(in == 313) begin
					state<=12;
					out<=37;
				end
				if(in == 314) begin
					state<=12;
					out<=38;
				end
				if(in == 315) begin
					state<=12;
					out<=39;
				end
				if(in == 316) begin
					state<=12;
					out<=40;
				end
				if(in == 317) begin
					state<=12;
					out<=41;
				end
				if(in == 318) begin
					state<=12;
					out<=42;
				end
				if(in == 319) begin
					state<=12;
					out<=43;
				end
				if(in == 320) begin
					state<=12;
					out<=44;
				end
				if(in == 321) begin
					state<=12;
					out<=45;
				end
				if(in == 322) begin
					state<=12;
					out<=46;
				end
				if(in == 323) begin
					state<=12;
					out<=47;
				end
				if(in == 324) begin
					state<=12;
					out<=48;
				end
				if(in == 325) begin
					state<=12;
					out<=49;
				end
				if(in == 326) begin
					state<=12;
					out<=50;
				end
				if(in == 327) begin
					state<=12;
					out<=51;
				end
				if(in == 328) begin
					state<=12;
					out<=52;
				end
				if(in == 329) begin
					state<=12;
					out<=53;
				end
				if(in == 330) begin
					state<=12;
					out<=54;
				end
				if(in == 331) begin
					state<=12;
					out<=55;
				end
				if(in == 332) begin
					state<=12;
					out<=56;
				end
				if(in == 333) begin
					state<=12;
					out<=57;
				end
				if(in == 334) begin
					state<=12;
					out<=58;
				end
				if(in == 335) begin
					state<=12;
					out<=59;
				end
				if(in == 336) begin
					state<=12;
					out<=60;
				end
				if(in == 337) begin
					state<=2;
					out<=61;
				end
				if(in == 338) begin
					state<=2;
					out<=62;
				end
				if(in == 339) begin
					state<=2;
					out<=63;
				end
				if(in == 340) begin
					state<=2;
					out<=64;
				end
				if(in == 341) begin
					state<=2;
					out<=65;
				end
				if(in == 342) begin
					state<=2;
					out<=66;
				end
				if(in == 343) begin
					state<=2;
					out<=67;
				end
				if(in == 344) begin
					state<=2;
					out<=68;
				end
				if(in == 345) begin
					state<=2;
					out<=69;
				end
				if(in == 346) begin
					state<=2;
					out<=70;
				end
				if(in == 347) begin
					state<=2;
					out<=71;
				end
				if(in == 348) begin
					state<=2;
					out<=72;
				end
				if(in == 349) begin
					state<=13;
					out<=73;
				end
				if(in == 350) begin
					state<=12;
					out<=74;
				end
				if(in == 351) begin
					state<=13;
					out<=75;
				end
				if(in == 352) begin
					state<=12;
					out<=76;
				end
				if(in == 353) begin
					state<=13;
					out<=77;
				end
				if(in == 354) begin
					state<=12;
					out<=78;
				end
				if(in == 355) begin
					state<=12;
					out<=79;
				end
				if(in == 356) begin
					state<=12;
					out<=80;
				end
				if(in == 357) begin
					state<=12;
					out<=81;
				end
				if(in == 358) begin
					state<=12;
					out<=82;
				end
				if(in == 359) begin
					state<=12;
					out<=83;
				end
				if(in == 360) begin
					state<=12;
					out<=84;
				end
				if(in == 361) begin
					state<=12;
					out<=85;
				end
				if(in == 362) begin
					state<=12;
					out<=86;
				end
				if(in == 363) begin
					state<=12;
					out<=87;
				end
				if(in == 364) begin
					state<=12;
					out<=88;
				end
				if(in == 365) begin
					state<=12;
					out<=89;
				end
				if(in == 366) begin
					state<=12;
					out<=90;
				end
				if(in == 367) begin
					state<=12;
					out<=91;
				end
				if(in == 368) begin
					state<=12;
					out<=92;
				end
				if(in == 369) begin
					state<=12;
					out<=93;
				end
				if(in == 370) begin
					state<=12;
					out<=94;
				end
				if(in == 371) begin
					state<=12;
					out<=95;
				end
				if(in == 372) begin
					state<=12;
					out<=96;
				end
				if(in == 373) begin
					state<=12;
					out<=97;
				end
				if(in == 374) begin
					state<=12;
					out<=98;
				end
				if(in == 375) begin
					state<=12;
					out<=99;
				end
				if(in == 376) begin
					state<=12;
					out<=100;
				end
				if(in == 377) begin
					state<=12;
					out<=101;
				end
				if(in == 378) begin
					state<=12;
					out<=102;
				end
				if(in == 379) begin
					state<=12;
					out<=103;
				end
				if(in == 380) begin
					state<=12;
					out<=104;
				end
				if(in == 381) begin
					state<=12;
					out<=105;
				end
				if(in == 382) begin
					state<=12;
					out<=106;
				end
				if(in == 383) begin
					state<=12;
					out<=107;
				end
				if(in == 384) begin
					state<=12;
					out<=108;
				end
				if(in == 385) begin
					state<=12;
					out<=109;
				end
				if(in == 386) begin
					state<=12;
					out<=110;
				end
				if(in == 387) begin
					state<=12;
					out<=111;
				end
				if(in == 388) begin
					state<=12;
					out<=112;
				end
				if(in == 389) begin
					state<=12;
					out<=113;
				end
				if(in == 390) begin
					state<=12;
					out<=114;
				end
				if(in == 391) begin
					state<=12;
					out<=115;
				end
				if(in == 392) begin
					state<=12;
					out<=116;
				end
				if(in == 393) begin
					state<=12;
					out<=117;
				end
				if(in == 394) begin
					state<=12;
					out<=118;
				end
				if(in == 395) begin
					state<=12;
					out<=119;
				end
				if(in == 396) begin
					state<=12;
					out<=120;
				end
				if(in == 397) begin
					state<=12;
					out<=121;
				end
				if(in == 398) begin
					state<=12;
					out<=122;
				end
				if(in == 399) begin
					state<=12;
					out<=123;
				end
				if(in == 400) begin
					state<=12;
					out<=124;
				end
				if(in == 401) begin
					state<=13;
					out<=125;
				end
				if(in == 402) begin
					state<=12;
					out<=126;
				end
				if(in == 403) begin
					state<=13;
					out<=127;
				end
				if(in == 404) begin
					state<=12;
					out<=128;
				end
				if(in == 405) begin
					state<=13;
					out<=129;
				end
				if(in == 406) begin
					state<=12;
					out<=130;
				end
				if(in == 407) begin
					state<=12;
					out<=131;
				end
				if(in == 408) begin
					state<=12;
					out<=132;
				end
				if(in == 409) begin
					state<=12;
					out<=133;
				end
				if(in == 410) begin
					state<=12;
					out<=134;
				end
				if(in == 411) begin
					state<=12;
					out<=135;
				end
				if(in == 412) begin
					state<=12;
					out<=136;
				end
				if(in == 413) begin
					state<=12;
					out<=137;
				end
				if(in == 414) begin
					state<=12;
					out<=138;
				end
				if(in == 415) begin
					state<=12;
					out<=139;
				end
				if(in == 416) begin
					state<=12;
					out<=140;
				end
				if(in == 417) begin
					state<=12;
					out<=141;
				end
				if(in == 418) begin
					state<=12;
					out<=142;
				end
				if(in == 419) begin
					state<=12;
					out<=143;
				end
				if(in == 420) begin
					state<=12;
					out<=144;
				end
				if(in == 421) begin
					state<=12;
					out<=145;
				end
				if(in == 422) begin
					state<=12;
					out<=146;
				end
				if(in == 423) begin
					state<=12;
					out<=147;
				end
				if(in == 424) begin
					state<=12;
					out<=148;
				end
				if(in == 425) begin
					state<=12;
					out<=149;
				end
				if(in == 426) begin
					state<=12;
					out<=150;
				end
				if(in == 427) begin
					state<=12;
					out<=151;
				end
				if(in == 428) begin
					state<=12;
					out<=152;
				end
				if(in == 429) begin
					state<=12;
					out<=153;
				end
				if(in == 430) begin
					state<=12;
					out<=154;
				end
				if(in == 431) begin
					state<=12;
					out<=155;
				end
				if(in == 432) begin
					state<=12;
					out<=156;
				end
				if(in == 433) begin
					state<=12;
					out<=157;
				end
				if(in == 434) begin
					state<=12;
					out<=158;
				end
				if(in == 435) begin
					state<=12;
					out<=159;
				end
				if(in == 436) begin
					state<=12;
					out<=160;
				end
				if(in == 437) begin
					state<=12;
					out<=161;
				end
				if(in == 438) begin
					state<=12;
					out<=162;
				end
				if(in == 439) begin
					state<=12;
					out<=163;
				end
				if(in == 440) begin
					state<=12;
					out<=164;
				end
				if(in == 441) begin
					state<=12;
					out<=165;
				end
				if(in == 442) begin
					state<=12;
					out<=166;
				end
				if(in == 443) begin
					state<=12;
					out<=167;
				end
				if(in == 444) begin
					state<=12;
					out<=168;
				end
				if(in == 445) begin
					state<=12;
					out<=169;
				end
				if(in == 446) begin
					state<=12;
					out<=170;
				end
				if(in == 447) begin
					state<=12;
					out<=171;
				end
				if(in == 448) begin
					state<=12;
					out<=172;
				end
				if(in == 449) begin
					state<=12;
					out<=173;
				end
				if(in == 450) begin
					state<=12;
					out<=174;
				end
				if(in == 451) begin
					state<=12;
					out<=175;
				end
				if(in == 452) begin
					state<=12;
					out<=176;
				end
				if(in == 453) begin
					state<=2;
					out<=177;
				end
				if(in == 454) begin
					state<=2;
					out<=178;
				end
				if(in == 455) begin
					state<=2;
					out<=179;
				end
				if(in == 456) begin
					state<=2;
					out<=180;
				end
				if(in == 457) begin
					state<=2;
					out<=181;
				end
				if(in == 458) begin
					state<=2;
					out<=182;
				end
				if(in == 459) begin
					state<=2;
					out<=183;
				end
				if(in == 460) begin
					state<=2;
					out<=184;
				end
				if(in == 461) begin
					state<=2;
					out<=185;
				end
				if(in == 462) begin
					state<=2;
					out<=186;
				end
				if(in == 463) begin
					state<=2;
					out<=187;
				end
				if(in == 464) begin
					state<=2;
					out<=188;
				end
				if(in == 465) begin
					state<=13;
					out<=189;
				end
				if(in == 466) begin
					state<=12;
					out<=190;
				end
				if(in == 467) begin
					state<=13;
					out<=191;
				end
				if(in == 468) begin
					state<=12;
					out<=192;
				end
				if(in == 469) begin
					state<=13;
					out<=193;
				end
				if(in == 470) begin
					state<=12;
					out<=194;
				end
				if(in == 471) begin
					state<=12;
					out<=195;
				end
				if(in == 472) begin
					state<=12;
					out<=196;
				end
				if(in == 473) begin
					state<=12;
					out<=197;
				end
				if(in == 474) begin
					state<=12;
					out<=198;
				end
				if(in == 475) begin
					state<=12;
					out<=199;
				end
				if(in == 476) begin
					state<=12;
					out<=200;
				end
				if(in == 477) begin
					state<=12;
					out<=201;
				end
				if(in == 478) begin
					state<=12;
					out<=202;
				end
				if(in == 479) begin
					state<=12;
					out<=203;
				end
				if(in == 480) begin
					state<=12;
					out<=204;
				end
				if(in == 481) begin
					state<=12;
					out<=205;
				end
				if(in == 482) begin
					state<=12;
					out<=206;
				end
				if(in == 483) begin
					state<=12;
					out<=207;
				end
				if(in == 484) begin
					state<=12;
					out<=208;
				end
				if(in == 485) begin
					state<=12;
					out<=209;
				end
				if(in == 486) begin
					state<=12;
					out<=210;
				end
				if(in == 487) begin
					state<=12;
					out<=211;
				end
				if(in == 488) begin
					state<=12;
					out<=212;
				end
				if(in == 489) begin
					state<=12;
					out<=213;
				end
				if(in == 490) begin
					state<=12;
					out<=214;
				end
				if(in == 491) begin
					state<=12;
					out<=215;
				end
				if(in == 492) begin
					state<=12;
					out<=216;
				end
				if(in == 493) begin
					state<=12;
					out<=217;
				end
				if(in == 494) begin
					state<=12;
					out<=218;
				end
				if(in == 495) begin
					state<=12;
					out<=219;
				end
				if(in == 496) begin
					state<=12;
					out<=220;
				end
				if(in == 497) begin
					state<=12;
					out<=221;
				end
				if(in == 498) begin
					state<=12;
					out<=222;
				end
				if(in == 499) begin
					state<=12;
					out<=223;
				end
				if(in == 500) begin
					state<=12;
					out<=224;
				end
				if(in == 501) begin
					state<=12;
					out<=225;
				end
				if(in == 502) begin
					state<=12;
					out<=226;
				end
				if(in == 503) begin
					state<=12;
					out<=227;
				end
				if(in == 504) begin
					state<=12;
					out<=228;
				end
				if(in == 505) begin
					state<=12;
					out<=229;
				end
				if(in == 506) begin
					state<=12;
					out<=230;
				end
				if(in == 507) begin
					state<=12;
					out<=231;
				end
				if(in == 508) begin
					state<=12;
					out<=232;
				end
				if(in == 509) begin
					state<=12;
					out<=233;
				end
				if(in == 510) begin
					state<=12;
					out<=234;
				end
				if(in == 511) begin
					state<=12;
					out<=235;
				end
				if(in == 512) begin
					state<=12;
					out<=236;
				end
				if(in == 513) begin
					state<=12;
					out<=237;
				end
				if(in == 514) begin
					state<=12;
					out<=238;
				end
				if(in == 515) begin
					state<=12;
					out<=239;
				end
				if(in == 516) begin
					state<=12;
					out<=240;
				end
				if(in == 517) begin
					state<=13;
					out<=241;
				end
				if(in == 518) begin
					state<=12;
					out<=242;
				end
				if(in == 519) begin
					state<=13;
					out<=243;
				end
				if(in == 520) begin
					state<=12;
					out<=244;
				end
				if(in == 521) begin
					state<=13;
					out<=245;
				end
				if(in == 522) begin
					state<=12;
					out<=246;
				end
				if(in == 523) begin
					state<=12;
					out<=247;
				end
				if(in == 524) begin
					state<=12;
					out<=248;
				end
				if(in == 525) begin
					state<=12;
					out<=249;
				end
				if(in == 526) begin
					state<=12;
					out<=250;
				end
				if(in == 527) begin
					state<=12;
					out<=251;
				end
				if(in == 528) begin
					state<=12;
					out<=252;
				end
				if(in == 529) begin
					state<=12;
					out<=253;
				end
				if(in == 530) begin
					state<=12;
					out<=254;
				end
				if(in == 531) begin
					state<=12;
					out<=255;
				end
				if(in == 532) begin
					state<=12;
					out<=0;
				end
				if(in == 533) begin
					state<=12;
					out<=1;
				end
				if(in == 534) begin
					state<=12;
					out<=2;
				end
				if(in == 535) begin
					state<=12;
					out<=3;
				end
				if(in == 536) begin
					state<=12;
					out<=4;
				end
				if(in == 537) begin
					state<=12;
					out<=5;
				end
				if(in == 538) begin
					state<=12;
					out<=6;
				end
				if(in == 539) begin
					state<=12;
					out<=7;
				end
				if(in == 540) begin
					state<=12;
					out<=8;
				end
				if(in == 541) begin
					state<=12;
					out<=9;
				end
				if(in == 542) begin
					state<=12;
					out<=10;
				end
				if(in == 543) begin
					state<=12;
					out<=11;
				end
				if(in == 544) begin
					state<=12;
					out<=12;
				end
				if(in == 545) begin
					state<=12;
					out<=13;
				end
				if(in == 546) begin
					state<=12;
					out<=14;
				end
				if(in == 547) begin
					state<=12;
					out<=15;
				end
				if(in == 548) begin
					state<=12;
					out<=16;
				end
				if(in == 549) begin
					state<=12;
					out<=17;
				end
				if(in == 550) begin
					state<=12;
					out<=18;
				end
				if(in == 551) begin
					state<=12;
					out<=19;
				end
				if(in == 552) begin
					state<=12;
					out<=20;
				end
				if(in == 553) begin
					state<=12;
					out<=21;
				end
				if(in == 554) begin
					state<=12;
					out<=22;
				end
				if(in == 555) begin
					state<=12;
					out<=23;
				end
				if(in == 556) begin
					state<=12;
					out<=24;
				end
				if(in == 557) begin
					state<=12;
					out<=25;
				end
				if(in == 558) begin
					state<=12;
					out<=26;
				end
				if(in == 559) begin
					state<=12;
					out<=27;
				end
				if(in == 560) begin
					state<=12;
					out<=28;
				end
				if(in == 561) begin
					state<=12;
					out<=29;
				end
				if(in == 562) begin
					state<=12;
					out<=30;
				end
				if(in == 563) begin
					state<=12;
					out<=31;
				end
				if(in == 564) begin
					state<=12;
					out<=32;
				end
				if(in == 565) begin
					state<=12;
					out<=33;
				end
				if(in == 566) begin
					state<=12;
					out<=34;
				end
				if(in == 567) begin
					state<=12;
					out<=35;
				end
				if(in == 568) begin
					state<=12;
					out<=36;
				end
				if(in == 569) begin
					state<=2;
					out<=37;
				end
				if(in == 570) begin
					state<=2;
					out<=38;
				end
				if(in == 571) begin
					state<=2;
					out<=39;
				end
				if(in == 572) begin
					state<=2;
					out<=40;
				end
				if(in == 573) begin
					state<=2;
					out<=41;
				end
				if(in == 574) begin
					state<=2;
					out<=42;
				end
				if(in == 575) begin
					state<=2;
					out<=43;
				end
				if(in == 576) begin
					state<=2;
					out<=44;
				end
				if(in == 577) begin
					state<=2;
					out<=45;
				end
				if(in == 578) begin
					state<=2;
					out<=46;
				end
				if(in == 579) begin
					state<=2;
					out<=47;
				end
				if(in == 580) begin
					state<=2;
					out<=48;
				end
				if(in == 581) begin
					state<=13;
					out<=49;
				end
				if(in == 582) begin
					state<=12;
					out<=50;
				end
				if(in == 583) begin
					state<=13;
					out<=51;
				end
				if(in == 584) begin
					state<=12;
					out<=52;
				end
				if(in == 585) begin
					state<=13;
					out<=53;
				end
				if(in == 586) begin
					state<=12;
					out<=54;
				end
				if(in == 587) begin
					state<=12;
					out<=55;
				end
				if(in == 588) begin
					state<=12;
					out<=56;
				end
				if(in == 589) begin
					state<=12;
					out<=57;
				end
				if(in == 590) begin
					state<=12;
					out<=58;
				end
				if(in == 591) begin
					state<=12;
					out<=59;
				end
				if(in == 592) begin
					state<=12;
					out<=60;
				end
				if(in == 593) begin
					state<=12;
					out<=61;
				end
				if(in == 594) begin
					state<=12;
					out<=62;
				end
				if(in == 595) begin
					state<=12;
					out<=63;
				end
				if(in == 596) begin
					state<=12;
					out<=64;
				end
				if(in == 597) begin
					state<=12;
					out<=65;
				end
				if(in == 598) begin
					state<=12;
					out<=66;
				end
				if(in == 599) begin
					state<=12;
					out<=67;
				end
				if(in == 600) begin
					state<=12;
					out<=68;
				end
				if(in == 601) begin
					state<=12;
					out<=69;
				end
				if(in == 602) begin
					state<=12;
					out<=70;
				end
				if(in == 603) begin
					state<=12;
					out<=71;
				end
				if(in == 604) begin
					state<=12;
					out<=72;
				end
				if(in == 605) begin
					state<=12;
					out<=73;
				end
				if(in == 606) begin
					state<=12;
					out<=74;
				end
				if(in == 607) begin
					state<=12;
					out<=75;
				end
				if(in == 608) begin
					state<=12;
					out<=76;
				end
				if(in == 609) begin
					state<=12;
					out<=77;
				end
				if(in == 610) begin
					state<=12;
					out<=78;
				end
				if(in == 611) begin
					state<=12;
					out<=79;
				end
				if(in == 612) begin
					state<=12;
					out<=80;
				end
				if(in == 613) begin
					state<=12;
					out<=81;
				end
				if(in == 614) begin
					state<=12;
					out<=82;
				end
				if(in == 615) begin
					state<=12;
					out<=83;
				end
				if(in == 616) begin
					state<=12;
					out<=84;
				end
				if(in == 617) begin
					state<=12;
					out<=85;
				end
				if(in == 618) begin
					state<=12;
					out<=86;
				end
				if(in == 619) begin
					state<=12;
					out<=87;
				end
				if(in == 620) begin
					state<=12;
					out<=88;
				end
				if(in == 621) begin
					state<=12;
					out<=89;
				end
				if(in == 622) begin
					state<=12;
					out<=90;
				end
				if(in == 623) begin
					state<=12;
					out<=91;
				end
				if(in == 624) begin
					state<=12;
					out<=92;
				end
				if(in == 625) begin
					state<=12;
					out<=93;
				end
				if(in == 626) begin
					state<=12;
					out<=94;
				end
				if(in == 627) begin
					state<=12;
					out<=95;
				end
				if(in == 628) begin
					state<=12;
					out<=96;
				end
				if(in == 629) begin
					state<=12;
					out<=97;
				end
				if(in == 630) begin
					state<=12;
					out<=98;
				end
				if(in == 631) begin
					state<=12;
					out<=99;
				end
				if(in == 632) begin
					state<=12;
					out<=100;
				end
				if(in == 633) begin
					state<=13;
					out<=101;
				end
				if(in == 634) begin
					state<=12;
					out<=102;
				end
				if(in == 635) begin
					state<=13;
					out<=103;
				end
				if(in == 636) begin
					state<=12;
					out<=104;
				end
				if(in == 637) begin
					state<=13;
					out<=105;
				end
				if(in == 638) begin
					state<=12;
					out<=106;
				end
				if(in == 639) begin
					state<=12;
					out<=107;
				end
				if(in == 640) begin
					state<=12;
					out<=108;
				end
				if(in == 641) begin
					state<=12;
					out<=109;
				end
				if(in == 642) begin
					state<=12;
					out<=110;
				end
				if(in == 643) begin
					state<=12;
					out<=111;
				end
				if(in == 644) begin
					state<=12;
					out<=112;
				end
				if(in == 645) begin
					state<=12;
					out<=113;
				end
				if(in == 646) begin
					state<=12;
					out<=114;
				end
				if(in == 647) begin
					state<=12;
					out<=115;
				end
				if(in == 648) begin
					state<=12;
					out<=116;
				end
				if(in == 649) begin
					state<=12;
					out<=117;
				end
				if(in == 650) begin
					state<=12;
					out<=118;
				end
				if(in == 651) begin
					state<=12;
					out<=119;
				end
				if(in == 652) begin
					state<=12;
					out<=120;
				end
				if(in == 653) begin
					state<=12;
					out<=121;
				end
				if(in == 654) begin
					state<=12;
					out<=122;
				end
				if(in == 655) begin
					state<=12;
					out<=123;
				end
				if(in == 656) begin
					state<=12;
					out<=124;
				end
				if(in == 657) begin
					state<=12;
					out<=125;
				end
				if(in == 658) begin
					state<=12;
					out<=126;
				end
				if(in == 659) begin
					state<=12;
					out<=127;
				end
				if(in == 660) begin
					state<=12;
					out<=128;
				end
				if(in == 661) begin
					state<=12;
					out<=129;
				end
				if(in == 662) begin
					state<=12;
					out<=130;
				end
				if(in == 663) begin
					state<=12;
					out<=131;
				end
				if(in == 664) begin
					state<=12;
					out<=132;
				end
				if(in == 665) begin
					state<=12;
					out<=133;
				end
				if(in == 666) begin
					state<=12;
					out<=134;
				end
				if(in == 667) begin
					state<=12;
					out<=135;
				end
				if(in == 668) begin
					state<=12;
					out<=136;
				end
				if(in == 669) begin
					state<=12;
					out<=137;
				end
				if(in == 670) begin
					state<=12;
					out<=138;
				end
				if(in == 671) begin
					state<=12;
					out<=139;
				end
				if(in == 672) begin
					state<=12;
					out<=140;
				end
				if(in == 673) begin
					state<=12;
					out<=141;
				end
				if(in == 674) begin
					state<=12;
					out<=142;
				end
				if(in == 675) begin
					state<=12;
					out<=143;
				end
				if(in == 676) begin
					state<=12;
					out<=144;
				end
				if(in == 677) begin
					state<=12;
					out<=145;
				end
				if(in == 678) begin
					state<=12;
					out<=146;
				end
				if(in == 679) begin
					state<=12;
					out<=147;
				end
				if(in == 680) begin
					state<=12;
					out<=148;
				end
				if(in == 681) begin
					state<=12;
					out<=149;
				end
				if(in == 682) begin
					state<=12;
					out<=150;
				end
				if(in == 683) begin
					state<=12;
					out<=151;
				end
				if(in == 684) begin
					state<=12;
					out<=152;
				end
				if(in == 685) begin
					state<=2;
					out<=153;
				end
				if(in == 686) begin
					state<=2;
					out<=154;
				end
				if(in == 687) begin
					state<=2;
					out<=155;
				end
				if(in == 688) begin
					state<=2;
					out<=156;
				end
				if(in == 689) begin
					state<=2;
					out<=157;
				end
				if(in == 690) begin
					state<=2;
					out<=158;
				end
				if(in == 691) begin
					state<=2;
					out<=159;
				end
				if(in == 692) begin
					state<=2;
					out<=160;
				end
				if(in == 693) begin
					state<=2;
					out<=161;
				end
				if(in == 694) begin
					state<=2;
					out<=162;
				end
				if(in == 695) begin
					state<=2;
					out<=163;
				end
				if(in == 696) begin
					state<=2;
					out<=164;
				end
				if(in == 697) begin
					state<=13;
					out<=165;
				end
				if(in == 698) begin
					state<=12;
					out<=166;
				end
				if(in == 699) begin
					state<=13;
					out<=167;
				end
				if(in == 700) begin
					state<=12;
					out<=168;
				end
				if(in == 701) begin
					state<=13;
					out<=169;
				end
				if(in == 702) begin
					state<=12;
					out<=170;
				end
				if(in == 703) begin
					state<=12;
					out<=171;
				end
				if(in == 704) begin
					state<=12;
					out<=172;
				end
				if(in == 705) begin
					state<=12;
					out<=173;
				end
				if(in == 706) begin
					state<=12;
					out<=174;
				end
				if(in == 707) begin
					state<=12;
					out<=175;
				end
				if(in == 708) begin
					state<=12;
					out<=176;
				end
				if(in == 709) begin
					state<=12;
					out<=177;
				end
				if(in == 710) begin
					state<=12;
					out<=178;
				end
				if(in == 711) begin
					state<=12;
					out<=179;
				end
				if(in == 712) begin
					state<=12;
					out<=180;
				end
				if(in == 713) begin
					state<=12;
					out<=181;
				end
				if(in == 714) begin
					state<=12;
					out<=182;
				end
				if(in == 715) begin
					state<=12;
					out<=183;
				end
				if(in == 716) begin
					state<=12;
					out<=184;
				end
				if(in == 717) begin
					state<=12;
					out<=185;
				end
				if(in == 718) begin
					state<=12;
					out<=186;
				end
				if(in == 719) begin
					state<=12;
					out<=187;
				end
				if(in == 720) begin
					state<=12;
					out<=188;
				end
				if(in == 721) begin
					state<=12;
					out<=189;
				end
				if(in == 722) begin
					state<=12;
					out<=190;
				end
				if(in == 723) begin
					state<=12;
					out<=191;
				end
				if(in == 724) begin
					state<=12;
					out<=192;
				end
				if(in == 725) begin
					state<=12;
					out<=193;
				end
				if(in == 726) begin
					state<=12;
					out<=194;
				end
				if(in == 727) begin
					state<=12;
					out<=195;
				end
				if(in == 728) begin
					state<=12;
					out<=196;
				end
				if(in == 729) begin
					state<=12;
					out<=197;
				end
				if(in == 730) begin
					state<=12;
					out<=198;
				end
				if(in == 731) begin
					state<=12;
					out<=199;
				end
				if(in == 732) begin
					state<=12;
					out<=200;
				end
				if(in == 733) begin
					state<=12;
					out<=201;
				end
				if(in == 734) begin
					state<=12;
					out<=202;
				end
				if(in == 735) begin
					state<=12;
					out<=203;
				end
				if(in == 736) begin
					state<=12;
					out<=204;
				end
				if(in == 737) begin
					state<=12;
					out<=205;
				end
				if(in == 738) begin
					state<=12;
					out<=206;
				end
				if(in == 739) begin
					state<=12;
					out<=207;
				end
				if(in == 740) begin
					state<=12;
					out<=208;
				end
				if(in == 741) begin
					state<=12;
					out<=209;
				end
				if(in == 742) begin
					state<=12;
					out<=210;
				end
				if(in == 743) begin
					state<=12;
					out<=211;
				end
				if(in == 744) begin
					state<=12;
					out<=212;
				end
				if(in == 745) begin
					state<=12;
					out<=213;
				end
				if(in == 746) begin
					state<=12;
					out<=214;
				end
				if(in == 747) begin
					state<=12;
					out<=215;
				end
				if(in == 748) begin
					state<=12;
					out<=216;
				end
				if(in == 749) begin
					state<=13;
					out<=217;
				end
				if(in == 750) begin
					state<=12;
					out<=218;
				end
				if(in == 751) begin
					state<=13;
					out<=219;
				end
				if(in == 752) begin
					state<=12;
					out<=220;
				end
				if(in == 753) begin
					state<=13;
					out<=221;
				end
				if(in == 754) begin
					state<=12;
					out<=222;
				end
				if(in == 755) begin
					state<=12;
					out<=223;
				end
				if(in == 756) begin
					state<=12;
					out<=224;
				end
				if(in == 757) begin
					state<=12;
					out<=225;
				end
				if(in == 758) begin
					state<=12;
					out<=226;
				end
				if(in == 759) begin
					state<=12;
					out<=227;
				end
				if(in == 760) begin
					state<=12;
					out<=228;
				end
				if(in == 761) begin
					state<=12;
					out<=229;
				end
				if(in == 762) begin
					state<=12;
					out<=230;
				end
				if(in == 763) begin
					state<=12;
					out<=231;
				end
				if(in == 764) begin
					state<=12;
					out<=232;
				end
				if(in == 765) begin
					state<=12;
					out<=233;
				end
				if(in == 766) begin
					state<=12;
					out<=234;
				end
				if(in == 767) begin
					state<=12;
					out<=235;
				end
				if(in == 768) begin
					state<=12;
					out<=236;
				end
				if(in == 769) begin
					state<=12;
					out<=237;
				end
				if(in == 770) begin
					state<=12;
					out<=238;
				end
				if(in == 771) begin
					state<=12;
					out<=239;
				end
				if(in == 772) begin
					state<=12;
					out<=240;
				end
				if(in == 773) begin
					state<=12;
					out<=241;
				end
				if(in == 774) begin
					state<=12;
					out<=242;
				end
				if(in == 775) begin
					state<=12;
					out<=243;
				end
				if(in == 776) begin
					state<=12;
					out<=244;
				end
				if(in == 777) begin
					state<=12;
					out<=245;
				end
				if(in == 778) begin
					state<=12;
					out<=246;
				end
				if(in == 779) begin
					state<=12;
					out<=247;
				end
				if(in == 780) begin
					state<=12;
					out<=248;
				end
				if(in == 781) begin
					state<=12;
					out<=249;
				end
				if(in == 782) begin
					state<=12;
					out<=250;
				end
				if(in == 783) begin
					state<=12;
					out<=251;
				end
				if(in == 784) begin
					state<=12;
					out<=252;
				end
				if(in == 785) begin
					state<=12;
					out<=253;
				end
				if(in == 786) begin
					state<=12;
					out<=254;
				end
				if(in == 787) begin
					state<=12;
					out<=255;
				end
				if(in == 788) begin
					state<=12;
					out<=0;
				end
				if(in == 789) begin
					state<=12;
					out<=1;
				end
				if(in == 790) begin
					state<=12;
					out<=2;
				end
				if(in == 791) begin
					state<=12;
					out<=3;
				end
				if(in == 792) begin
					state<=12;
					out<=4;
				end
				if(in == 793) begin
					state<=12;
					out<=5;
				end
				if(in == 794) begin
					state<=12;
					out<=6;
				end
				if(in == 795) begin
					state<=12;
					out<=7;
				end
				if(in == 796) begin
					state<=12;
					out<=8;
				end
				if(in == 797) begin
					state<=12;
					out<=9;
				end
				if(in == 798) begin
					state<=12;
					out<=10;
				end
				if(in == 799) begin
					state<=12;
					out<=11;
				end
				if(in == 800) begin
					state<=12;
					out<=12;
				end
				if(in == 801) begin
					state<=2;
					out<=13;
				end
				if(in == 802) begin
					state<=2;
					out<=14;
				end
				if(in == 803) begin
					state<=2;
					out<=15;
				end
				if(in == 804) begin
					state<=2;
					out<=16;
				end
				if(in == 805) begin
					state<=2;
					out<=17;
				end
				if(in == 806) begin
					state<=2;
					out<=18;
				end
				if(in == 807) begin
					state<=2;
					out<=19;
				end
				if(in == 808) begin
					state<=2;
					out<=20;
				end
				if(in == 809) begin
					state<=2;
					out<=21;
				end
				if(in == 810) begin
					state<=2;
					out<=22;
				end
				if(in == 811) begin
					state<=2;
					out<=23;
				end
				if(in == 812) begin
					state<=2;
					out<=24;
				end
				if(in == 813) begin
					state<=13;
					out<=25;
				end
				if(in == 814) begin
					state<=12;
					out<=26;
				end
				if(in == 815) begin
					state<=13;
					out<=27;
				end
				if(in == 816) begin
					state<=12;
					out<=28;
				end
				if(in == 817) begin
					state<=13;
					out<=29;
				end
				if(in == 818) begin
					state<=12;
					out<=30;
				end
				if(in == 819) begin
					state<=12;
					out<=31;
				end
				if(in == 820) begin
					state<=12;
					out<=32;
				end
				if(in == 821) begin
					state<=12;
					out<=33;
				end
				if(in == 822) begin
					state<=12;
					out<=34;
				end
				if(in == 823) begin
					state<=12;
					out<=35;
				end
				if(in == 824) begin
					state<=12;
					out<=36;
				end
				if(in == 825) begin
					state<=12;
					out<=37;
				end
				if(in == 826) begin
					state<=12;
					out<=38;
				end
				if(in == 827) begin
					state<=12;
					out<=39;
				end
				if(in == 828) begin
					state<=12;
					out<=40;
				end
				if(in == 829) begin
					state<=12;
					out<=41;
				end
				if(in == 830) begin
					state<=12;
					out<=42;
				end
				if(in == 831) begin
					state<=12;
					out<=43;
				end
				if(in == 832) begin
					state<=12;
					out<=44;
				end
				if(in == 833) begin
					state<=12;
					out<=45;
				end
				if(in == 834) begin
					state<=12;
					out<=46;
				end
				if(in == 835) begin
					state<=12;
					out<=47;
				end
				if(in == 836) begin
					state<=12;
					out<=48;
				end
				if(in == 837) begin
					state<=12;
					out<=49;
				end
				if(in == 838) begin
					state<=12;
					out<=50;
				end
				if(in == 839) begin
					state<=12;
					out<=51;
				end
				if(in == 840) begin
					state<=12;
					out<=52;
				end
				if(in == 841) begin
					state<=12;
					out<=53;
				end
				if(in == 842) begin
					state<=12;
					out<=54;
				end
				if(in == 843) begin
					state<=12;
					out<=55;
				end
				if(in == 844) begin
					state<=12;
					out<=56;
				end
				if(in == 845) begin
					state<=12;
					out<=57;
				end
				if(in == 846) begin
					state<=12;
					out<=58;
				end
				if(in == 847) begin
					state<=12;
					out<=59;
				end
				if(in == 848) begin
					state<=12;
					out<=60;
				end
				if(in == 849) begin
					state<=12;
					out<=61;
				end
				if(in == 850) begin
					state<=12;
					out<=62;
				end
				if(in == 851) begin
					state<=12;
					out<=63;
				end
				if(in == 852) begin
					state<=12;
					out<=64;
				end
				if(in == 853) begin
					state<=12;
					out<=65;
				end
				if(in == 854) begin
					state<=12;
					out<=66;
				end
				if(in == 855) begin
					state<=12;
					out<=67;
				end
				if(in == 856) begin
					state<=12;
					out<=68;
				end
				if(in == 857) begin
					state<=12;
					out<=69;
				end
				if(in == 858) begin
					state<=12;
					out<=70;
				end
				if(in == 859) begin
					state<=12;
					out<=71;
				end
				if(in == 860) begin
					state<=12;
					out<=72;
				end
				if(in == 861) begin
					state<=12;
					out<=73;
				end
				if(in == 862) begin
					state<=12;
					out<=74;
				end
				if(in == 863) begin
					state<=12;
					out<=75;
				end
				if(in == 864) begin
					state<=12;
					out<=76;
				end
				if(in == 865) begin
					state<=13;
					out<=77;
				end
				if(in == 866) begin
					state<=12;
					out<=78;
				end
				if(in == 867) begin
					state<=13;
					out<=79;
				end
				if(in == 868) begin
					state<=12;
					out<=80;
				end
				if(in == 869) begin
					state<=13;
					out<=81;
				end
				if(in == 870) begin
					state<=12;
					out<=82;
				end
				if(in == 871) begin
					state<=12;
					out<=83;
				end
				if(in == 872) begin
					state<=12;
					out<=84;
				end
				if(in == 873) begin
					state<=12;
					out<=85;
				end
				if(in == 874) begin
					state<=12;
					out<=86;
				end
				if(in == 875) begin
					state<=12;
					out<=87;
				end
				if(in == 876) begin
					state<=12;
					out<=88;
				end
				if(in == 877) begin
					state<=12;
					out<=89;
				end
				if(in == 878) begin
					state<=12;
					out<=90;
				end
				if(in == 879) begin
					state<=12;
					out<=91;
				end
				if(in == 880) begin
					state<=12;
					out<=92;
				end
				if(in == 881) begin
					state<=12;
					out<=93;
				end
				if(in == 882) begin
					state<=12;
					out<=94;
				end
				if(in == 883) begin
					state<=12;
					out<=95;
				end
				if(in == 884) begin
					state<=12;
					out<=96;
				end
				if(in == 885) begin
					state<=12;
					out<=97;
				end
				if(in == 886) begin
					state<=12;
					out<=98;
				end
				if(in == 887) begin
					state<=12;
					out<=99;
				end
				if(in == 888) begin
					state<=12;
					out<=100;
				end
				if(in == 889) begin
					state<=12;
					out<=101;
				end
				if(in == 890) begin
					state<=12;
					out<=102;
				end
				if(in == 891) begin
					state<=12;
					out<=103;
				end
				if(in == 892) begin
					state<=12;
					out<=104;
				end
				if(in == 893) begin
					state<=12;
					out<=105;
				end
				if(in == 894) begin
					state<=12;
					out<=106;
				end
				if(in == 895) begin
					state<=12;
					out<=107;
				end
				if(in == 896) begin
					state<=12;
					out<=108;
				end
				if(in == 897) begin
					state<=12;
					out<=109;
				end
				if(in == 898) begin
					state<=12;
					out<=110;
				end
				if(in == 899) begin
					state<=12;
					out<=111;
				end
				if(in == 900) begin
					state<=12;
					out<=112;
				end
				if(in == 901) begin
					state<=12;
					out<=113;
				end
				if(in == 902) begin
					state<=12;
					out<=114;
				end
				if(in == 903) begin
					state<=12;
					out<=115;
				end
				if(in == 904) begin
					state<=12;
					out<=116;
				end
				if(in == 905) begin
					state<=12;
					out<=117;
				end
				if(in == 906) begin
					state<=12;
					out<=118;
				end
				if(in == 907) begin
					state<=12;
					out<=119;
				end
				if(in == 908) begin
					state<=12;
					out<=120;
				end
				if(in == 909) begin
					state<=12;
					out<=121;
				end
				if(in == 910) begin
					state<=12;
					out<=122;
				end
				if(in == 911) begin
					state<=12;
					out<=123;
				end
				if(in == 912) begin
					state<=12;
					out<=124;
				end
				if(in == 913) begin
					state<=12;
					out<=125;
				end
				if(in == 914) begin
					state<=12;
					out<=126;
				end
				if(in == 915) begin
					state<=12;
					out<=127;
				end
				if(in == 916) begin
					state<=12;
					out<=128;
				end
				if(in == 917) begin
					state<=2;
					out<=129;
				end
				if(in == 918) begin
					state<=2;
					out<=130;
				end
				if(in == 919) begin
					state<=2;
					out<=131;
				end
				if(in == 920) begin
					state<=2;
					out<=132;
				end
				if(in == 921) begin
					state<=2;
					out<=133;
				end
				if(in == 922) begin
					state<=2;
					out<=134;
				end
				if(in == 923) begin
					state<=2;
					out<=135;
				end
				if(in == 924) begin
					state<=2;
					out<=136;
				end
				if(in == 925) begin
					state<=2;
					out<=137;
				end
				if(in == 926) begin
					state<=2;
					out<=138;
				end
				if(in == 927) begin
					state<=2;
					out<=139;
				end
				if(in == 928) begin
					state<=2;
					out<=140;
				end
			end
			13: begin
				if(in == 0) begin
					state<=14;
					out<=141;
				end
				if(in == 1) begin
					state<=1;
					out<=142;
				end
				if(in == 2) begin
					state<=14;
					out<=143;
				end
				if(in == 3) begin
					state<=14;
					out<=144;
				end
				if(in == 4) begin
					state<=14;
					out<=145;
				end
				if(in == 5) begin
					state<=14;
					out<=146;
				end
				if(in == 6) begin
					state<=14;
					out<=147;
				end
				if(in == 7) begin
					state<=14;
					out<=148;
				end
				if(in == 8) begin
					state<=14;
					out<=149;
				end
				if(in == 9) begin
					state<=14;
					out<=150;
				end
				if(in == 10) begin
					state<=14;
					out<=151;
				end
				if(in == 11) begin
					state<=14;
					out<=152;
				end
				if(in == 12) begin
					state<=14;
					out<=153;
				end
				if(in == 13) begin
					state<=14;
					out<=154;
				end
				if(in == 14) begin
					state<=14;
					out<=155;
				end
				if(in == 15) begin
					state<=14;
					out<=156;
				end
				if(in == 16) begin
					state<=14;
					out<=157;
				end
				if(in == 17) begin
					state<=14;
					out<=158;
				end
				if(in == 18) begin
					state<=14;
					out<=159;
				end
				if(in == 19) begin
					state<=14;
					out<=160;
				end
				if(in == 20) begin
					state<=14;
					out<=161;
				end
				if(in == 21) begin
					state<=14;
					out<=162;
				end
				if(in == 22) begin
					state<=14;
					out<=163;
				end
				if(in == 23) begin
					state<=14;
					out<=164;
				end
				if(in == 24) begin
					state<=14;
					out<=165;
				end
				if(in == 25) begin
					state<=14;
					out<=166;
				end
				if(in == 26) begin
					state<=14;
					out<=167;
				end
				if(in == 27) begin
					state<=14;
					out<=168;
				end
				if(in == 28) begin
					state<=14;
					out<=169;
				end
				if(in == 29) begin
					state<=14;
					out<=170;
				end
				if(in == 30) begin
					state<=14;
					out<=171;
				end
				if(in == 31) begin
					state<=14;
					out<=172;
				end
				if(in == 32) begin
					state<=14;
					out<=173;
				end
				if(in == 33) begin
					state<=14;
					out<=174;
				end
				if(in == 34) begin
					state<=14;
					out<=175;
				end
				if(in == 35) begin
					state<=14;
					out<=176;
				end
				if(in == 36) begin
					state<=14;
					out<=177;
				end
				if(in == 37) begin
					state<=14;
					out<=178;
				end
				if(in == 38) begin
					state<=14;
					out<=179;
				end
				if(in == 39) begin
					state<=14;
					out<=180;
				end
				if(in == 40) begin
					state<=14;
					out<=181;
				end
				if(in == 41) begin
					state<=14;
					out<=182;
				end
				if(in == 42) begin
					state<=14;
					out<=183;
				end
				if(in == 43) begin
					state<=14;
					out<=184;
				end
				if(in == 44) begin
					state<=14;
					out<=185;
				end
				if(in == 45) begin
					state<=14;
					out<=186;
				end
				if(in == 46) begin
					state<=14;
					out<=187;
				end
				if(in == 47) begin
					state<=14;
					out<=188;
				end
				if(in == 48) begin
					state<=14;
					out<=189;
				end
				if(in == 49) begin
					state<=14;
					out<=190;
				end
				if(in == 50) begin
					state<=14;
					out<=191;
				end
				if(in == 51) begin
					state<=14;
					out<=192;
				end
				if(in == 52) begin
					state<=14;
					out<=193;
				end
				if(in == 53) begin
					state<=3;
					out<=194;
				end
				if(in == 54) begin
					state<=3;
					out<=195;
				end
				if(in == 55) begin
					state<=3;
					out<=196;
				end
				if(in == 56) begin
					state<=3;
					out<=197;
				end
				if(in == 57) begin
					state<=3;
					out<=198;
				end
				if(in == 58) begin
					state<=3;
					out<=199;
				end
				if(in == 59) begin
					state<=3;
					out<=200;
				end
				if(in == 60) begin
					state<=3;
					out<=201;
				end
				if(in == 61) begin
					state<=3;
					out<=202;
				end
				if(in == 62) begin
					state<=3;
					out<=203;
				end
				if(in == 63) begin
					state<=3;
					out<=204;
				end
				if(in == 64) begin
					state<=3;
					out<=205;
				end
				if(in == 65) begin
					state<=3;
					out<=206;
				end
				if(in == 66) begin
					state<=3;
					out<=207;
				end
				if(in == 67) begin
					state<=3;
					out<=208;
				end
				if(in == 68) begin
					state<=3;
					out<=209;
				end
				if(in == 69) begin
					state<=3;
					out<=210;
				end
				if(in == 70) begin
					state<=3;
					out<=211;
				end
				if(in == 71) begin
					state<=3;
					out<=212;
				end
				if(in == 72) begin
					state<=3;
					out<=213;
				end
				if(in == 73) begin
					state<=3;
					out<=214;
				end
				if(in == 74) begin
					state<=3;
					out<=215;
				end
				if(in == 75) begin
					state<=3;
					out<=216;
				end
				if(in == 76) begin
					state<=3;
					out<=217;
				end
				if(in == 77) begin
					state<=3;
					out<=218;
				end
				if(in == 78) begin
					state<=3;
					out<=219;
				end
				if(in == 79) begin
					state<=3;
					out<=220;
				end
				if(in == 80) begin
					state<=3;
					out<=221;
				end
				if(in == 81) begin
					state<=3;
					out<=222;
				end
				if(in == 82) begin
					state<=3;
					out<=223;
				end
				if(in == 83) begin
					state<=3;
					out<=224;
				end
				if(in == 84) begin
					state<=3;
					out<=225;
				end
				if(in == 85) begin
					state<=3;
					out<=226;
				end
				if(in == 86) begin
					state<=3;
					out<=227;
				end
				if(in == 87) begin
					state<=3;
					out<=228;
				end
				if(in == 88) begin
					state<=3;
					out<=229;
				end
				if(in == 89) begin
					state<=3;
					out<=230;
				end
				if(in == 90) begin
					state<=3;
					out<=231;
				end
				if(in == 91) begin
					state<=3;
					out<=232;
				end
				if(in == 92) begin
					state<=3;
					out<=233;
				end
				if(in == 93) begin
					state<=3;
					out<=234;
				end
				if(in == 94) begin
					state<=3;
					out<=235;
				end
				if(in == 95) begin
					state<=3;
					out<=236;
				end
				if(in == 96) begin
					state<=3;
					out<=237;
				end
				if(in == 97) begin
					state<=3;
					out<=238;
				end
				if(in == 98) begin
					state<=3;
					out<=239;
				end
				if(in == 99) begin
					state<=3;
					out<=240;
				end
				if(in == 100) begin
					state<=3;
					out<=241;
				end
				if(in == 101) begin
					state<=3;
					out<=242;
				end
				if(in == 102) begin
					state<=3;
					out<=243;
				end
				if(in == 103) begin
					state<=3;
					out<=244;
				end
				if(in == 104) begin
					state<=3;
					out<=245;
				end
				if(in == 105) begin
					state<=14;
					out<=246;
				end
				if(in == 106) begin
					state<=14;
					out<=247;
				end
				if(in == 107) begin
					state<=14;
					out<=248;
				end
				if(in == 108) begin
					state<=14;
					out<=249;
				end
				if(in == 109) begin
					state<=14;
					out<=250;
				end
				if(in == 110) begin
					state<=14;
					out<=251;
				end
				if(in == 111) begin
					state<=3;
					out<=252;
				end
				if(in == 112) begin
					state<=3;
					out<=253;
				end
				if(in == 113) begin
					state<=3;
					out<=254;
				end
				if(in == 114) begin
					state<=3;
					out<=255;
				end
				if(in == 115) begin
					state<=3;
					out<=0;
				end
				if(in == 116) begin
					state<=3;
					out<=1;
				end
				if(in == 117) begin
					state<=14;
					out<=2;
				end
				if(in == 118) begin
					state<=14;
					out<=3;
				end
				if(in == 119) begin
					state<=14;
					out<=4;
				end
				if(in == 120) begin
					state<=14;
					out<=5;
				end
				if(in == 121) begin
					state<=14;
					out<=6;
				end
				if(in == 122) begin
					state<=14;
					out<=7;
				end
				if(in == 123) begin
					state<=14;
					out<=8;
				end
				if(in == 124) begin
					state<=14;
					out<=9;
				end
				if(in == 125) begin
					state<=14;
					out<=10;
				end
				if(in == 126) begin
					state<=14;
					out<=11;
				end
				if(in == 127) begin
					state<=14;
					out<=12;
				end
				if(in == 128) begin
					state<=14;
					out<=13;
				end
				if(in == 129) begin
					state<=14;
					out<=14;
				end
				if(in == 130) begin
					state<=14;
					out<=15;
				end
				if(in == 131) begin
					state<=14;
					out<=16;
				end
				if(in == 132) begin
					state<=14;
					out<=17;
				end
				if(in == 133) begin
					state<=14;
					out<=18;
				end
				if(in == 134) begin
					state<=14;
					out<=19;
				end
				if(in == 135) begin
					state<=14;
					out<=20;
				end
				if(in == 136) begin
					state<=14;
					out<=21;
				end
				if(in == 137) begin
					state<=14;
					out<=22;
				end
				if(in == 138) begin
					state<=14;
					out<=23;
				end
				if(in == 139) begin
					state<=14;
					out<=24;
				end
				if(in == 140) begin
					state<=14;
					out<=25;
				end
				if(in == 141) begin
					state<=14;
					out<=26;
				end
				if(in == 142) begin
					state<=14;
					out<=27;
				end
				if(in == 143) begin
					state<=14;
					out<=28;
				end
				if(in == 144) begin
					state<=14;
					out<=29;
				end
				if(in == 145) begin
					state<=14;
					out<=30;
				end
				if(in == 146) begin
					state<=14;
					out<=31;
				end
				if(in == 147) begin
					state<=14;
					out<=32;
				end
				if(in == 148) begin
					state<=14;
					out<=33;
				end
				if(in == 149) begin
					state<=14;
					out<=34;
				end
				if(in == 150) begin
					state<=14;
					out<=35;
				end
				if(in == 151) begin
					state<=14;
					out<=36;
				end
				if(in == 152) begin
					state<=14;
					out<=37;
				end
				if(in == 153) begin
					state<=14;
					out<=38;
				end
				if(in == 154) begin
					state<=14;
					out<=39;
				end
				if(in == 155) begin
					state<=14;
					out<=40;
				end
				if(in == 156) begin
					state<=14;
					out<=41;
				end
				if(in == 157) begin
					state<=14;
					out<=42;
				end
				if(in == 158) begin
					state<=14;
					out<=43;
				end
				if(in == 159) begin
					state<=14;
					out<=44;
				end
				if(in == 160) begin
					state<=14;
					out<=45;
				end
				if(in == 161) begin
					state<=14;
					out<=46;
				end
				if(in == 162) begin
					state<=14;
					out<=47;
				end
				if(in == 163) begin
					state<=14;
					out<=48;
				end
				if(in == 164) begin
					state<=14;
					out<=49;
				end
				if(in == 165) begin
					state<=14;
					out<=50;
				end
				if(in == 166) begin
					state<=14;
					out<=51;
				end
				if(in == 167) begin
					state<=14;
					out<=52;
				end
				if(in == 168) begin
					state<=14;
					out<=53;
				end
				if(in == 169) begin
					state<=3;
					out<=54;
				end
				if(in == 170) begin
					state<=3;
					out<=55;
				end
				if(in == 171) begin
					state<=3;
					out<=56;
				end
				if(in == 172) begin
					state<=3;
					out<=57;
				end
				if(in == 173) begin
					state<=3;
					out<=58;
				end
				if(in == 174) begin
					state<=3;
					out<=59;
				end
				if(in == 175) begin
					state<=3;
					out<=60;
				end
				if(in == 176) begin
					state<=3;
					out<=61;
				end
				if(in == 177) begin
					state<=3;
					out<=62;
				end
				if(in == 178) begin
					state<=3;
					out<=63;
				end
				if(in == 179) begin
					state<=3;
					out<=64;
				end
				if(in == 180) begin
					state<=3;
					out<=65;
				end
				if(in == 181) begin
					state<=3;
					out<=66;
				end
				if(in == 182) begin
					state<=3;
					out<=67;
				end
				if(in == 183) begin
					state<=3;
					out<=68;
				end
				if(in == 184) begin
					state<=3;
					out<=69;
				end
				if(in == 185) begin
					state<=3;
					out<=70;
				end
				if(in == 186) begin
					state<=3;
					out<=71;
				end
				if(in == 187) begin
					state<=3;
					out<=72;
				end
				if(in == 188) begin
					state<=3;
					out<=73;
				end
				if(in == 189) begin
					state<=3;
					out<=74;
				end
				if(in == 190) begin
					state<=3;
					out<=75;
				end
				if(in == 191) begin
					state<=3;
					out<=76;
				end
				if(in == 192) begin
					state<=3;
					out<=77;
				end
				if(in == 193) begin
					state<=3;
					out<=78;
				end
				if(in == 194) begin
					state<=3;
					out<=79;
				end
				if(in == 195) begin
					state<=3;
					out<=80;
				end
				if(in == 196) begin
					state<=3;
					out<=81;
				end
				if(in == 197) begin
					state<=3;
					out<=82;
				end
				if(in == 198) begin
					state<=3;
					out<=83;
				end
				if(in == 199) begin
					state<=3;
					out<=84;
				end
				if(in == 200) begin
					state<=3;
					out<=85;
				end
				if(in == 201) begin
					state<=3;
					out<=86;
				end
				if(in == 202) begin
					state<=3;
					out<=87;
				end
				if(in == 203) begin
					state<=3;
					out<=88;
				end
				if(in == 204) begin
					state<=3;
					out<=89;
				end
				if(in == 205) begin
					state<=3;
					out<=90;
				end
				if(in == 206) begin
					state<=3;
					out<=91;
				end
				if(in == 207) begin
					state<=3;
					out<=92;
				end
				if(in == 208) begin
					state<=3;
					out<=93;
				end
				if(in == 209) begin
					state<=3;
					out<=94;
				end
				if(in == 210) begin
					state<=3;
					out<=95;
				end
				if(in == 211) begin
					state<=3;
					out<=96;
				end
				if(in == 212) begin
					state<=3;
					out<=97;
				end
				if(in == 213) begin
					state<=3;
					out<=98;
				end
				if(in == 214) begin
					state<=3;
					out<=99;
				end
				if(in == 215) begin
					state<=3;
					out<=100;
				end
				if(in == 216) begin
					state<=3;
					out<=101;
				end
				if(in == 217) begin
					state<=3;
					out<=102;
				end
				if(in == 218) begin
					state<=3;
					out<=103;
				end
				if(in == 219) begin
					state<=3;
					out<=104;
				end
				if(in == 220) begin
					state<=3;
					out<=105;
				end
				if(in == 221) begin
					state<=14;
					out<=106;
				end
				if(in == 222) begin
					state<=14;
					out<=107;
				end
				if(in == 223) begin
					state<=14;
					out<=108;
				end
				if(in == 224) begin
					state<=14;
					out<=109;
				end
				if(in == 225) begin
					state<=14;
					out<=110;
				end
				if(in == 226) begin
					state<=14;
					out<=111;
				end
				if(in == 227) begin
					state<=3;
					out<=112;
				end
				if(in == 228) begin
					state<=3;
					out<=113;
				end
				if(in == 229) begin
					state<=3;
					out<=114;
				end
				if(in == 230) begin
					state<=3;
					out<=115;
				end
				if(in == 231) begin
					state<=3;
					out<=116;
				end
				if(in == 232) begin
					state<=3;
					out<=117;
				end
				if(in == 233) begin
					state<=14;
					out<=118;
				end
				if(in == 234) begin
					state<=14;
					out<=119;
				end
				if(in == 235) begin
					state<=14;
					out<=120;
				end
				if(in == 236) begin
					state<=14;
					out<=121;
				end
				if(in == 237) begin
					state<=14;
					out<=122;
				end
				if(in == 238) begin
					state<=14;
					out<=123;
				end
				if(in == 239) begin
					state<=14;
					out<=124;
				end
				if(in == 240) begin
					state<=14;
					out<=125;
				end
				if(in == 241) begin
					state<=14;
					out<=126;
				end
				if(in == 242) begin
					state<=14;
					out<=127;
				end
				if(in == 243) begin
					state<=14;
					out<=128;
				end
				if(in == 244) begin
					state<=14;
					out<=129;
				end
				if(in == 245) begin
					state<=14;
					out<=130;
				end
				if(in == 246) begin
					state<=14;
					out<=131;
				end
				if(in == 247) begin
					state<=14;
					out<=132;
				end
				if(in == 248) begin
					state<=14;
					out<=133;
				end
				if(in == 249) begin
					state<=14;
					out<=134;
				end
				if(in == 250) begin
					state<=14;
					out<=135;
				end
				if(in == 251) begin
					state<=14;
					out<=136;
				end
				if(in == 252) begin
					state<=14;
					out<=137;
				end
				if(in == 253) begin
					state<=14;
					out<=138;
				end
				if(in == 254) begin
					state<=14;
					out<=139;
				end
				if(in == 255) begin
					state<=14;
					out<=140;
				end
				if(in == 256) begin
					state<=14;
					out<=141;
				end
				if(in == 257) begin
					state<=14;
					out<=142;
				end
				if(in == 258) begin
					state<=14;
					out<=143;
				end
				if(in == 259) begin
					state<=14;
					out<=144;
				end
				if(in == 260) begin
					state<=14;
					out<=145;
				end
				if(in == 261) begin
					state<=14;
					out<=146;
				end
				if(in == 262) begin
					state<=14;
					out<=147;
				end
				if(in == 263) begin
					state<=14;
					out<=148;
				end
				if(in == 264) begin
					state<=14;
					out<=149;
				end
				if(in == 265) begin
					state<=14;
					out<=150;
				end
				if(in == 266) begin
					state<=14;
					out<=151;
				end
				if(in == 267) begin
					state<=14;
					out<=152;
				end
				if(in == 268) begin
					state<=14;
					out<=153;
				end
				if(in == 269) begin
					state<=14;
					out<=154;
				end
				if(in == 270) begin
					state<=14;
					out<=155;
				end
				if(in == 271) begin
					state<=14;
					out<=156;
				end
				if(in == 272) begin
					state<=14;
					out<=157;
				end
				if(in == 273) begin
					state<=14;
					out<=158;
				end
				if(in == 274) begin
					state<=14;
					out<=159;
				end
				if(in == 275) begin
					state<=14;
					out<=160;
				end
				if(in == 276) begin
					state<=14;
					out<=161;
				end
				if(in == 277) begin
					state<=14;
					out<=162;
				end
				if(in == 278) begin
					state<=14;
					out<=163;
				end
				if(in == 279) begin
					state<=14;
					out<=164;
				end
				if(in == 280) begin
					state<=14;
					out<=165;
				end
				if(in == 281) begin
					state<=14;
					out<=166;
				end
				if(in == 282) begin
					state<=14;
					out<=167;
				end
				if(in == 283) begin
					state<=14;
					out<=168;
				end
				if(in == 284) begin
					state<=14;
					out<=169;
				end
				if(in == 285) begin
					state<=3;
					out<=170;
				end
				if(in == 286) begin
					state<=3;
					out<=171;
				end
				if(in == 287) begin
					state<=3;
					out<=172;
				end
				if(in == 288) begin
					state<=3;
					out<=173;
				end
				if(in == 289) begin
					state<=3;
					out<=174;
				end
				if(in == 290) begin
					state<=3;
					out<=175;
				end
				if(in == 291) begin
					state<=3;
					out<=176;
				end
				if(in == 292) begin
					state<=3;
					out<=177;
				end
				if(in == 293) begin
					state<=3;
					out<=178;
				end
				if(in == 294) begin
					state<=3;
					out<=179;
				end
				if(in == 295) begin
					state<=3;
					out<=180;
				end
				if(in == 296) begin
					state<=3;
					out<=181;
				end
				if(in == 297) begin
					state<=3;
					out<=182;
				end
				if(in == 298) begin
					state<=3;
					out<=183;
				end
				if(in == 299) begin
					state<=3;
					out<=184;
				end
				if(in == 300) begin
					state<=3;
					out<=185;
				end
				if(in == 301) begin
					state<=3;
					out<=186;
				end
				if(in == 302) begin
					state<=3;
					out<=187;
				end
				if(in == 303) begin
					state<=3;
					out<=188;
				end
				if(in == 304) begin
					state<=3;
					out<=189;
				end
				if(in == 305) begin
					state<=3;
					out<=190;
				end
				if(in == 306) begin
					state<=3;
					out<=191;
				end
				if(in == 307) begin
					state<=3;
					out<=192;
				end
				if(in == 308) begin
					state<=3;
					out<=193;
				end
				if(in == 309) begin
					state<=3;
					out<=194;
				end
				if(in == 310) begin
					state<=3;
					out<=195;
				end
				if(in == 311) begin
					state<=3;
					out<=196;
				end
				if(in == 312) begin
					state<=3;
					out<=197;
				end
				if(in == 313) begin
					state<=3;
					out<=198;
				end
				if(in == 314) begin
					state<=3;
					out<=199;
				end
				if(in == 315) begin
					state<=3;
					out<=200;
				end
				if(in == 316) begin
					state<=3;
					out<=201;
				end
				if(in == 317) begin
					state<=3;
					out<=202;
				end
				if(in == 318) begin
					state<=3;
					out<=203;
				end
				if(in == 319) begin
					state<=3;
					out<=204;
				end
				if(in == 320) begin
					state<=3;
					out<=205;
				end
				if(in == 321) begin
					state<=3;
					out<=206;
				end
				if(in == 322) begin
					state<=3;
					out<=207;
				end
				if(in == 323) begin
					state<=3;
					out<=208;
				end
				if(in == 324) begin
					state<=3;
					out<=209;
				end
				if(in == 325) begin
					state<=3;
					out<=210;
				end
				if(in == 326) begin
					state<=3;
					out<=211;
				end
				if(in == 327) begin
					state<=3;
					out<=212;
				end
				if(in == 328) begin
					state<=3;
					out<=213;
				end
				if(in == 329) begin
					state<=3;
					out<=214;
				end
				if(in == 330) begin
					state<=3;
					out<=215;
				end
				if(in == 331) begin
					state<=3;
					out<=216;
				end
				if(in == 332) begin
					state<=3;
					out<=217;
				end
				if(in == 333) begin
					state<=3;
					out<=218;
				end
				if(in == 334) begin
					state<=3;
					out<=219;
				end
				if(in == 335) begin
					state<=3;
					out<=220;
				end
				if(in == 336) begin
					state<=3;
					out<=221;
				end
				if(in == 337) begin
					state<=14;
					out<=222;
				end
				if(in == 338) begin
					state<=14;
					out<=223;
				end
				if(in == 339) begin
					state<=14;
					out<=224;
				end
				if(in == 340) begin
					state<=14;
					out<=225;
				end
				if(in == 341) begin
					state<=14;
					out<=226;
				end
				if(in == 342) begin
					state<=14;
					out<=227;
				end
				if(in == 343) begin
					state<=3;
					out<=228;
				end
				if(in == 344) begin
					state<=3;
					out<=229;
				end
				if(in == 345) begin
					state<=3;
					out<=230;
				end
				if(in == 346) begin
					state<=3;
					out<=231;
				end
				if(in == 347) begin
					state<=3;
					out<=232;
				end
				if(in == 348) begin
					state<=3;
					out<=233;
				end
				if(in == 349) begin
					state<=14;
					out<=234;
				end
				if(in == 350) begin
					state<=14;
					out<=235;
				end
				if(in == 351) begin
					state<=14;
					out<=236;
				end
				if(in == 352) begin
					state<=14;
					out<=237;
				end
				if(in == 353) begin
					state<=14;
					out<=238;
				end
				if(in == 354) begin
					state<=14;
					out<=239;
				end
				if(in == 355) begin
					state<=14;
					out<=240;
				end
				if(in == 356) begin
					state<=14;
					out<=241;
				end
				if(in == 357) begin
					state<=14;
					out<=242;
				end
				if(in == 358) begin
					state<=14;
					out<=243;
				end
				if(in == 359) begin
					state<=14;
					out<=244;
				end
				if(in == 360) begin
					state<=14;
					out<=245;
				end
				if(in == 361) begin
					state<=14;
					out<=246;
				end
				if(in == 362) begin
					state<=14;
					out<=247;
				end
				if(in == 363) begin
					state<=14;
					out<=248;
				end
				if(in == 364) begin
					state<=14;
					out<=249;
				end
				if(in == 365) begin
					state<=14;
					out<=250;
				end
				if(in == 366) begin
					state<=14;
					out<=251;
				end
				if(in == 367) begin
					state<=14;
					out<=252;
				end
				if(in == 368) begin
					state<=14;
					out<=253;
				end
				if(in == 369) begin
					state<=14;
					out<=254;
				end
				if(in == 370) begin
					state<=14;
					out<=255;
				end
				if(in == 371) begin
					state<=14;
					out<=0;
				end
				if(in == 372) begin
					state<=14;
					out<=1;
				end
				if(in == 373) begin
					state<=14;
					out<=2;
				end
				if(in == 374) begin
					state<=14;
					out<=3;
				end
				if(in == 375) begin
					state<=14;
					out<=4;
				end
				if(in == 376) begin
					state<=14;
					out<=5;
				end
				if(in == 377) begin
					state<=14;
					out<=6;
				end
				if(in == 378) begin
					state<=14;
					out<=7;
				end
				if(in == 379) begin
					state<=14;
					out<=8;
				end
				if(in == 380) begin
					state<=14;
					out<=9;
				end
				if(in == 381) begin
					state<=14;
					out<=10;
				end
				if(in == 382) begin
					state<=14;
					out<=11;
				end
				if(in == 383) begin
					state<=14;
					out<=12;
				end
				if(in == 384) begin
					state<=14;
					out<=13;
				end
				if(in == 385) begin
					state<=14;
					out<=14;
				end
				if(in == 386) begin
					state<=14;
					out<=15;
				end
				if(in == 387) begin
					state<=14;
					out<=16;
				end
				if(in == 388) begin
					state<=14;
					out<=17;
				end
				if(in == 389) begin
					state<=14;
					out<=18;
				end
				if(in == 390) begin
					state<=14;
					out<=19;
				end
				if(in == 391) begin
					state<=14;
					out<=20;
				end
				if(in == 392) begin
					state<=14;
					out<=21;
				end
				if(in == 393) begin
					state<=14;
					out<=22;
				end
				if(in == 394) begin
					state<=14;
					out<=23;
				end
				if(in == 395) begin
					state<=14;
					out<=24;
				end
				if(in == 396) begin
					state<=14;
					out<=25;
				end
				if(in == 397) begin
					state<=14;
					out<=26;
				end
				if(in == 398) begin
					state<=14;
					out<=27;
				end
				if(in == 399) begin
					state<=14;
					out<=28;
				end
				if(in == 400) begin
					state<=14;
					out<=29;
				end
				if(in == 401) begin
					state<=3;
					out<=30;
				end
				if(in == 402) begin
					state<=3;
					out<=31;
				end
				if(in == 403) begin
					state<=3;
					out<=32;
				end
				if(in == 404) begin
					state<=3;
					out<=33;
				end
				if(in == 405) begin
					state<=3;
					out<=34;
				end
				if(in == 406) begin
					state<=3;
					out<=35;
				end
				if(in == 407) begin
					state<=3;
					out<=36;
				end
				if(in == 408) begin
					state<=3;
					out<=37;
				end
				if(in == 409) begin
					state<=3;
					out<=38;
				end
				if(in == 410) begin
					state<=3;
					out<=39;
				end
				if(in == 411) begin
					state<=3;
					out<=40;
				end
				if(in == 412) begin
					state<=3;
					out<=41;
				end
				if(in == 413) begin
					state<=3;
					out<=42;
				end
				if(in == 414) begin
					state<=3;
					out<=43;
				end
				if(in == 415) begin
					state<=3;
					out<=44;
				end
				if(in == 416) begin
					state<=3;
					out<=45;
				end
				if(in == 417) begin
					state<=3;
					out<=46;
				end
				if(in == 418) begin
					state<=3;
					out<=47;
				end
				if(in == 419) begin
					state<=3;
					out<=48;
				end
				if(in == 420) begin
					state<=3;
					out<=49;
				end
				if(in == 421) begin
					state<=3;
					out<=50;
				end
				if(in == 422) begin
					state<=3;
					out<=51;
				end
				if(in == 423) begin
					state<=3;
					out<=52;
				end
				if(in == 424) begin
					state<=3;
					out<=53;
				end
				if(in == 425) begin
					state<=3;
					out<=54;
				end
				if(in == 426) begin
					state<=3;
					out<=55;
				end
				if(in == 427) begin
					state<=3;
					out<=56;
				end
				if(in == 428) begin
					state<=3;
					out<=57;
				end
				if(in == 429) begin
					state<=3;
					out<=58;
				end
				if(in == 430) begin
					state<=3;
					out<=59;
				end
				if(in == 431) begin
					state<=3;
					out<=60;
				end
				if(in == 432) begin
					state<=3;
					out<=61;
				end
				if(in == 433) begin
					state<=3;
					out<=62;
				end
				if(in == 434) begin
					state<=3;
					out<=63;
				end
				if(in == 435) begin
					state<=3;
					out<=64;
				end
				if(in == 436) begin
					state<=3;
					out<=65;
				end
				if(in == 437) begin
					state<=3;
					out<=66;
				end
				if(in == 438) begin
					state<=3;
					out<=67;
				end
				if(in == 439) begin
					state<=3;
					out<=68;
				end
				if(in == 440) begin
					state<=3;
					out<=69;
				end
				if(in == 441) begin
					state<=3;
					out<=70;
				end
				if(in == 442) begin
					state<=3;
					out<=71;
				end
				if(in == 443) begin
					state<=3;
					out<=72;
				end
				if(in == 444) begin
					state<=3;
					out<=73;
				end
				if(in == 445) begin
					state<=3;
					out<=74;
				end
				if(in == 446) begin
					state<=3;
					out<=75;
				end
				if(in == 447) begin
					state<=3;
					out<=76;
				end
				if(in == 448) begin
					state<=3;
					out<=77;
				end
				if(in == 449) begin
					state<=3;
					out<=78;
				end
				if(in == 450) begin
					state<=3;
					out<=79;
				end
				if(in == 451) begin
					state<=3;
					out<=80;
				end
				if(in == 452) begin
					state<=3;
					out<=81;
				end
				if(in == 453) begin
					state<=14;
					out<=82;
				end
				if(in == 454) begin
					state<=14;
					out<=83;
				end
				if(in == 455) begin
					state<=14;
					out<=84;
				end
				if(in == 456) begin
					state<=14;
					out<=85;
				end
				if(in == 457) begin
					state<=14;
					out<=86;
				end
				if(in == 458) begin
					state<=14;
					out<=87;
				end
				if(in == 459) begin
					state<=3;
					out<=88;
				end
				if(in == 460) begin
					state<=3;
					out<=89;
				end
				if(in == 461) begin
					state<=3;
					out<=90;
				end
				if(in == 462) begin
					state<=3;
					out<=91;
				end
				if(in == 463) begin
					state<=3;
					out<=92;
				end
				if(in == 464) begin
					state<=3;
					out<=93;
				end
				if(in == 465) begin
					state<=14;
					out<=94;
				end
				if(in == 466) begin
					state<=14;
					out<=95;
				end
				if(in == 467) begin
					state<=14;
					out<=96;
				end
				if(in == 468) begin
					state<=14;
					out<=97;
				end
				if(in == 469) begin
					state<=14;
					out<=98;
				end
				if(in == 470) begin
					state<=14;
					out<=99;
				end
				if(in == 471) begin
					state<=14;
					out<=100;
				end
				if(in == 472) begin
					state<=14;
					out<=101;
				end
				if(in == 473) begin
					state<=14;
					out<=102;
				end
				if(in == 474) begin
					state<=14;
					out<=103;
				end
				if(in == 475) begin
					state<=14;
					out<=104;
				end
				if(in == 476) begin
					state<=14;
					out<=105;
				end
				if(in == 477) begin
					state<=14;
					out<=106;
				end
				if(in == 478) begin
					state<=14;
					out<=107;
				end
				if(in == 479) begin
					state<=14;
					out<=108;
				end
				if(in == 480) begin
					state<=14;
					out<=109;
				end
				if(in == 481) begin
					state<=14;
					out<=110;
				end
				if(in == 482) begin
					state<=14;
					out<=111;
				end
				if(in == 483) begin
					state<=14;
					out<=112;
				end
				if(in == 484) begin
					state<=14;
					out<=113;
				end
				if(in == 485) begin
					state<=14;
					out<=114;
				end
				if(in == 486) begin
					state<=14;
					out<=115;
				end
				if(in == 487) begin
					state<=14;
					out<=116;
				end
				if(in == 488) begin
					state<=14;
					out<=117;
				end
				if(in == 489) begin
					state<=14;
					out<=118;
				end
				if(in == 490) begin
					state<=14;
					out<=119;
				end
				if(in == 491) begin
					state<=14;
					out<=120;
				end
				if(in == 492) begin
					state<=14;
					out<=121;
				end
				if(in == 493) begin
					state<=14;
					out<=122;
				end
				if(in == 494) begin
					state<=14;
					out<=123;
				end
				if(in == 495) begin
					state<=14;
					out<=124;
				end
				if(in == 496) begin
					state<=14;
					out<=125;
				end
				if(in == 497) begin
					state<=14;
					out<=126;
				end
				if(in == 498) begin
					state<=14;
					out<=127;
				end
				if(in == 499) begin
					state<=14;
					out<=128;
				end
				if(in == 500) begin
					state<=14;
					out<=129;
				end
				if(in == 501) begin
					state<=14;
					out<=130;
				end
				if(in == 502) begin
					state<=14;
					out<=131;
				end
				if(in == 503) begin
					state<=14;
					out<=132;
				end
				if(in == 504) begin
					state<=14;
					out<=133;
				end
				if(in == 505) begin
					state<=14;
					out<=134;
				end
				if(in == 506) begin
					state<=14;
					out<=135;
				end
				if(in == 507) begin
					state<=14;
					out<=136;
				end
				if(in == 508) begin
					state<=14;
					out<=137;
				end
				if(in == 509) begin
					state<=14;
					out<=138;
				end
				if(in == 510) begin
					state<=14;
					out<=139;
				end
				if(in == 511) begin
					state<=14;
					out<=140;
				end
				if(in == 512) begin
					state<=14;
					out<=141;
				end
				if(in == 513) begin
					state<=14;
					out<=142;
				end
				if(in == 514) begin
					state<=14;
					out<=143;
				end
				if(in == 515) begin
					state<=14;
					out<=144;
				end
				if(in == 516) begin
					state<=14;
					out<=145;
				end
				if(in == 517) begin
					state<=3;
					out<=146;
				end
				if(in == 518) begin
					state<=3;
					out<=147;
				end
				if(in == 519) begin
					state<=3;
					out<=148;
				end
				if(in == 520) begin
					state<=3;
					out<=149;
				end
				if(in == 521) begin
					state<=3;
					out<=150;
				end
				if(in == 522) begin
					state<=3;
					out<=151;
				end
				if(in == 523) begin
					state<=3;
					out<=152;
				end
				if(in == 524) begin
					state<=3;
					out<=153;
				end
				if(in == 525) begin
					state<=3;
					out<=154;
				end
				if(in == 526) begin
					state<=3;
					out<=155;
				end
				if(in == 527) begin
					state<=3;
					out<=156;
				end
				if(in == 528) begin
					state<=3;
					out<=157;
				end
				if(in == 529) begin
					state<=3;
					out<=158;
				end
				if(in == 530) begin
					state<=3;
					out<=159;
				end
				if(in == 531) begin
					state<=3;
					out<=160;
				end
				if(in == 532) begin
					state<=3;
					out<=161;
				end
				if(in == 533) begin
					state<=3;
					out<=162;
				end
				if(in == 534) begin
					state<=3;
					out<=163;
				end
				if(in == 535) begin
					state<=3;
					out<=164;
				end
				if(in == 536) begin
					state<=3;
					out<=165;
				end
				if(in == 537) begin
					state<=3;
					out<=166;
				end
				if(in == 538) begin
					state<=3;
					out<=167;
				end
				if(in == 539) begin
					state<=3;
					out<=168;
				end
				if(in == 540) begin
					state<=3;
					out<=169;
				end
				if(in == 541) begin
					state<=3;
					out<=170;
				end
				if(in == 542) begin
					state<=3;
					out<=171;
				end
				if(in == 543) begin
					state<=3;
					out<=172;
				end
				if(in == 544) begin
					state<=3;
					out<=173;
				end
				if(in == 545) begin
					state<=3;
					out<=174;
				end
				if(in == 546) begin
					state<=3;
					out<=175;
				end
				if(in == 547) begin
					state<=3;
					out<=176;
				end
				if(in == 548) begin
					state<=3;
					out<=177;
				end
				if(in == 549) begin
					state<=3;
					out<=178;
				end
				if(in == 550) begin
					state<=3;
					out<=179;
				end
				if(in == 551) begin
					state<=3;
					out<=180;
				end
				if(in == 552) begin
					state<=3;
					out<=181;
				end
				if(in == 553) begin
					state<=3;
					out<=182;
				end
				if(in == 554) begin
					state<=3;
					out<=183;
				end
				if(in == 555) begin
					state<=3;
					out<=184;
				end
				if(in == 556) begin
					state<=3;
					out<=185;
				end
				if(in == 557) begin
					state<=3;
					out<=186;
				end
				if(in == 558) begin
					state<=3;
					out<=187;
				end
				if(in == 559) begin
					state<=3;
					out<=188;
				end
				if(in == 560) begin
					state<=3;
					out<=189;
				end
				if(in == 561) begin
					state<=3;
					out<=190;
				end
				if(in == 562) begin
					state<=3;
					out<=191;
				end
				if(in == 563) begin
					state<=3;
					out<=192;
				end
				if(in == 564) begin
					state<=3;
					out<=193;
				end
				if(in == 565) begin
					state<=3;
					out<=194;
				end
				if(in == 566) begin
					state<=3;
					out<=195;
				end
				if(in == 567) begin
					state<=3;
					out<=196;
				end
				if(in == 568) begin
					state<=3;
					out<=197;
				end
				if(in == 569) begin
					state<=14;
					out<=198;
				end
				if(in == 570) begin
					state<=14;
					out<=199;
				end
				if(in == 571) begin
					state<=14;
					out<=200;
				end
				if(in == 572) begin
					state<=14;
					out<=201;
				end
				if(in == 573) begin
					state<=14;
					out<=202;
				end
				if(in == 574) begin
					state<=14;
					out<=203;
				end
				if(in == 575) begin
					state<=3;
					out<=204;
				end
				if(in == 576) begin
					state<=3;
					out<=205;
				end
				if(in == 577) begin
					state<=3;
					out<=206;
				end
				if(in == 578) begin
					state<=3;
					out<=207;
				end
				if(in == 579) begin
					state<=3;
					out<=208;
				end
				if(in == 580) begin
					state<=3;
					out<=209;
				end
				if(in == 581) begin
					state<=14;
					out<=210;
				end
				if(in == 582) begin
					state<=14;
					out<=211;
				end
				if(in == 583) begin
					state<=14;
					out<=212;
				end
				if(in == 584) begin
					state<=14;
					out<=213;
				end
				if(in == 585) begin
					state<=14;
					out<=214;
				end
				if(in == 586) begin
					state<=14;
					out<=215;
				end
				if(in == 587) begin
					state<=14;
					out<=216;
				end
				if(in == 588) begin
					state<=14;
					out<=217;
				end
				if(in == 589) begin
					state<=14;
					out<=218;
				end
				if(in == 590) begin
					state<=14;
					out<=219;
				end
				if(in == 591) begin
					state<=14;
					out<=220;
				end
				if(in == 592) begin
					state<=14;
					out<=221;
				end
				if(in == 593) begin
					state<=14;
					out<=222;
				end
				if(in == 594) begin
					state<=14;
					out<=223;
				end
				if(in == 595) begin
					state<=14;
					out<=224;
				end
				if(in == 596) begin
					state<=14;
					out<=225;
				end
				if(in == 597) begin
					state<=14;
					out<=226;
				end
				if(in == 598) begin
					state<=14;
					out<=227;
				end
				if(in == 599) begin
					state<=14;
					out<=228;
				end
				if(in == 600) begin
					state<=14;
					out<=229;
				end
				if(in == 601) begin
					state<=14;
					out<=230;
				end
				if(in == 602) begin
					state<=14;
					out<=231;
				end
				if(in == 603) begin
					state<=14;
					out<=232;
				end
				if(in == 604) begin
					state<=14;
					out<=233;
				end
				if(in == 605) begin
					state<=14;
					out<=234;
				end
				if(in == 606) begin
					state<=14;
					out<=235;
				end
				if(in == 607) begin
					state<=14;
					out<=236;
				end
				if(in == 608) begin
					state<=14;
					out<=237;
				end
				if(in == 609) begin
					state<=14;
					out<=238;
				end
				if(in == 610) begin
					state<=14;
					out<=239;
				end
				if(in == 611) begin
					state<=14;
					out<=240;
				end
				if(in == 612) begin
					state<=14;
					out<=241;
				end
				if(in == 613) begin
					state<=14;
					out<=242;
				end
				if(in == 614) begin
					state<=14;
					out<=243;
				end
				if(in == 615) begin
					state<=14;
					out<=244;
				end
				if(in == 616) begin
					state<=14;
					out<=245;
				end
				if(in == 617) begin
					state<=14;
					out<=246;
				end
				if(in == 618) begin
					state<=14;
					out<=247;
				end
				if(in == 619) begin
					state<=14;
					out<=248;
				end
				if(in == 620) begin
					state<=14;
					out<=249;
				end
				if(in == 621) begin
					state<=14;
					out<=250;
				end
				if(in == 622) begin
					state<=14;
					out<=251;
				end
				if(in == 623) begin
					state<=14;
					out<=252;
				end
				if(in == 624) begin
					state<=14;
					out<=253;
				end
				if(in == 625) begin
					state<=14;
					out<=254;
				end
				if(in == 626) begin
					state<=14;
					out<=255;
				end
				if(in == 627) begin
					state<=14;
					out<=0;
				end
				if(in == 628) begin
					state<=14;
					out<=1;
				end
				if(in == 629) begin
					state<=14;
					out<=2;
				end
				if(in == 630) begin
					state<=14;
					out<=3;
				end
				if(in == 631) begin
					state<=14;
					out<=4;
				end
				if(in == 632) begin
					state<=14;
					out<=5;
				end
				if(in == 633) begin
					state<=3;
					out<=6;
				end
				if(in == 634) begin
					state<=3;
					out<=7;
				end
				if(in == 635) begin
					state<=3;
					out<=8;
				end
				if(in == 636) begin
					state<=3;
					out<=9;
				end
				if(in == 637) begin
					state<=3;
					out<=10;
				end
				if(in == 638) begin
					state<=3;
					out<=11;
				end
				if(in == 639) begin
					state<=3;
					out<=12;
				end
				if(in == 640) begin
					state<=3;
					out<=13;
				end
				if(in == 641) begin
					state<=3;
					out<=14;
				end
				if(in == 642) begin
					state<=3;
					out<=15;
				end
				if(in == 643) begin
					state<=3;
					out<=16;
				end
				if(in == 644) begin
					state<=3;
					out<=17;
				end
				if(in == 645) begin
					state<=3;
					out<=18;
				end
				if(in == 646) begin
					state<=3;
					out<=19;
				end
				if(in == 647) begin
					state<=3;
					out<=20;
				end
				if(in == 648) begin
					state<=3;
					out<=21;
				end
				if(in == 649) begin
					state<=3;
					out<=22;
				end
				if(in == 650) begin
					state<=3;
					out<=23;
				end
				if(in == 651) begin
					state<=3;
					out<=24;
				end
				if(in == 652) begin
					state<=3;
					out<=25;
				end
				if(in == 653) begin
					state<=3;
					out<=26;
				end
				if(in == 654) begin
					state<=3;
					out<=27;
				end
				if(in == 655) begin
					state<=3;
					out<=28;
				end
				if(in == 656) begin
					state<=3;
					out<=29;
				end
				if(in == 657) begin
					state<=3;
					out<=30;
				end
				if(in == 658) begin
					state<=3;
					out<=31;
				end
				if(in == 659) begin
					state<=3;
					out<=32;
				end
				if(in == 660) begin
					state<=3;
					out<=33;
				end
				if(in == 661) begin
					state<=3;
					out<=34;
				end
				if(in == 662) begin
					state<=3;
					out<=35;
				end
				if(in == 663) begin
					state<=3;
					out<=36;
				end
				if(in == 664) begin
					state<=3;
					out<=37;
				end
				if(in == 665) begin
					state<=3;
					out<=38;
				end
				if(in == 666) begin
					state<=3;
					out<=39;
				end
				if(in == 667) begin
					state<=3;
					out<=40;
				end
				if(in == 668) begin
					state<=3;
					out<=41;
				end
				if(in == 669) begin
					state<=3;
					out<=42;
				end
				if(in == 670) begin
					state<=3;
					out<=43;
				end
				if(in == 671) begin
					state<=3;
					out<=44;
				end
				if(in == 672) begin
					state<=3;
					out<=45;
				end
				if(in == 673) begin
					state<=3;
					out<=46;
				end
				if(in == 674) begin
					state<=3;
					out<=47;
				end
				if(in == 675) begin
					state<=3;
					out<=48;
				end
				if(in == 676) begin
					state<=3;
					out<=49;
				end
				if(in == 677) begin
					state<=3;
					out<=50;
				end
				if(in == 678) begin
					state<=3;
					out<=51;
				end
				if(in == 679) begin
					state<=3;
					out<=52;
				end
				if(in == 680) begin
					state<=3;
					out<=53;
				end
				if(in == 681) begin
					state<=3;
					out<=54;
				end
				if(in == 682) begin
					state<=3;
					out<=55;
				end
				if(in == 683) begin
					state<=3;
					out<=56;
				end
				if(in == 684) begin
					state<=3;
					out<=57;
				end
				if(in == 685) begin
					state<=14;
					out<=58;
				end
				if(in == 686) begin
					state<=14;
					out<=59;
				end
				if(in == 687) begin
					state<=14;
					out<=60;
				end
				if(in == 688) begin
					state<=14;
					out<=61;
				end
				if(in == 689) begin
					state<=14;
					out<=62;
				end
				if(in == 690) begin
					state<=14;
					out<=63;
				end
				if(in == 691) begin
					state<=3;
					out<=64;
				end
				if(in == 692) begin
					state<=3;
					out<=65;
				end
				if(in == 693) begin
					state<=3;
					out<=66;
				end
				if(in == 694) begin
					state<=3;
					out<=67;
				end
				if(in == 695) begin
					state<=3;
					out<=68;
				end
				if(in == 696) begin
					state<=3;
					out<=69;
				end
				if(in == 697) begin
					state<=14;
					out<=70;
				end
				if(in == 698) begin
					state<=14;
					out<=71;
				end
				if(in == 699) begin
					state<=14;
					out<=72;
				end
				if(in == 700) begin
					state<=14;
					out<=73;
				end
				if(in == 701) begin
					state<=14;
					out<=74;
				end
				if(in == 702) begin
					state<=14;
					out<=75;
				end
				if(in == 703) begin
					state<=14;
					out<=76;
				end
				if(in == 704) begin
					state<=14;
					out<=77;
				end
				if(in == 705) begin
					state<=14;
					out<=78;
				end
				if(in == 706) begin
					state<=14;
					out<=79;
				end
				if(in == 707) begin
					state<=14;
					out<=80;
				end
				if(in == 708) begin
					state<=14;
					out<=81;
				end
				if(in == 709) begin
					state<=14;
					out<=82;
				end
				if(in == 710) begin
					state<=14;
					out<=83;
				end
				if(in == 711) begin
					state<=14;
					out<=84;
				end
				if(in == 712) begin
					state<=14;
					out<=85;
				end
				if(in == 713) begin
					state<=14;
					out<=86;
				end
				if(in == 714) begin
					state<=14;
					out<=87;
				end
				if(in == 715) begin
					state<=14;
					out<=88;
				end
				if(in == 716) begin
					state<=14;
					out<=89;
				end
				if(in == 717) begin
					state<=14;
					out<=90;
				end
				if(in == 718) begin
					state<=14;
					out<=91;
				end
				if(in == 719) begin
					state<=14;
					out<=92;
				end
				if(in == 720) begin
					state<=14;
					out<=93;
				end
				if(in == 721) begin
					state<=14;
					out<=94;
				end
				if(in == 722) begin
					state<=14;
					out<=95;
				end
				if(in == 723) begin
					state<=14;
					out<=96;
				end
				if(in == 724) begin
					state<=14;
					out<=97;
				end
				if(in == 725) begin
					state<=14;
					out<=98;
				end
				if(in == 726) begin
					state<=14;
					out<=99;
				end
				if(in == 727) begin
					state<=14;
					out<=100;
				end
				if(in == 728) begin
					state<=14;
					out<=101;
				end
				if(in == 729) begin
					state<=14;
					out<=102;
				end
				if(in == 730) begin
					state<=14;
					out<=103;
				end
				if(in == 731) begin
					state<=14;
					out<=104;
				end
				if(in == 732) begin
					state<=14;
					out<=105;
				end
				if(in == 733) begin
					state<=14;
					out<=106;
				end
				if(in == 734) begin
					state<=14;
					out<=107;
				end
				if(in == 735) begin
					state<=14;
					out<=108;
				end
				if(in == 736) begin
					state<=14;
					out<=109;
				end
				if(in == 737) begin
					state<=14;
					out<=110;
				end
				if(in == 738) begin
					state<=14;
					out<=111;
				end
				if(in == 739) begin
					state<=14;
					out<=112;
				end
				if(in == 740) begin
					state<=14;
					out<=113;
				end
				if(in == 741) begin
					state<=14;
					out<=114;
				end
				if(in == 742) begin
					state<=14;
					out<=115;
				end
				if(in == 743) begin
					state<=14;
					out<=116;
				end
				if(in == 744) begin
					state<=14;
					out<=117;
				end
				if(in == 745) begin
					state<=14;
					out<=118;
				end
				if(in == 746) begin
					state<=14;
					out<=119;
				end
				if(in == 747) begin
					state<=14;
					out<=120;
				end
				if(in == 748) begin
					state<=14;
					out<=121;
				end
				if(in == 749) begin
					state<=3;
					out<=122;
				end
				if(in == 750) begin
					state<=3;
					out<=123;
				end
				if(in == 751) begin
					state<=3;
					out<=124;
				end
				if(in == 752) begin
					state<=3;
					out<=125;
				end
				if(in == 753) begin
					state<=3;
					out<=126;
				end
				if(in == 754) begin
					state<=3;
					out<=127;
				end
				if(in == 755) begin
					state<=3;
					out<=128;
				end
				if(in == 756) begin
					state<=3;
					out<=129;
				end
				if(in == 757) begin
					state<=3;
					out<=130;
				end
				if(in == 758) begin
					state<=3;
					out<=131;
				end
				if(in == 759) begin
					state<=3;
					out<=132;
				end
				if(in == 760) begin
					state<=3;
					out<=133;
				end
				if(in == 761) begin
					state<=3;
					out<=134;
				end
				if(in == 762) begin
					state<=3;
					out<=135;
				end
				if(in == 763) begin
					state<=3;
					out<=136;
				end
				if(in == 764) begin
					state<=3;
					out<=137;
				end
				if(in == 765) begin
					state<=3;
					out<=138;
				end
				if(in == 766) begin
					state<=3;
					out<=139;
				end
				if(in == 767) begin
					state<=3;
					out<=140;
				end
				if(in == 768) begin
					state<=3;
					out<=141;
				end
				if(in == 769) begin
					state<=3;
					out<=142;
				end
				if(in == 770) begin
					state<=3;
					out<=143;
				end
				if(in == 771) begin
					state<=3;
					out<=144;
				end
				if(in == 772) begin
					state<=3;
					out<=145;
				end
				if(in == 773) begin
					state<=3;
					out<=146;
				end
				if(in == 774) begin
					state<=3;
					out<=147;
				end
				if(in == 775) begin
					state<=3;
					out<=148;
				end
				if(in == 776) begin
					state<=3;
					out<=149;
				end
				if(in == 777) begin
					state<=3;
					out<=150;
				end
				if(in == 778) begin
					state<=3;
					out<=151;
				end
				if(in == 779) begin
					state<=3;
					out<=152;
				end
				if(in == 780) begin
					state<=3;
					out<=153;
				end
				if(in == 781) begin
					state<=3;
					out<=154;
				end
				if(in == 782) begin
					state<=3;
					out<=155;
				end
				if(in == 783) begin
					state<=3;
					out<=156;
				end
				if(in == 784) begin
					state<=3;
					out<=157;
				end
				if(in == 785) begin
					state<=3;
					out<=158;
				end
				if(in == 786) begin
					state<=3;
					out<=159;
				end
				if(in == 787) begin
					state<=3;
					out<=160;
				end
				if(in == 788) begin
					state<=3;
					out<=161;
				end
				if(in == 789) begin
					state<=3;
					out<=162;
				end
				if(in == 790) begin
					state<=3;
					out<=163;
				end
				if(in == 791) begin
					state<=3;
					out<=164;
				end
				if(in == 792) begin
					state<=3;
					out<=165;
				end
				if(in == 793) begin
					state<=3;
					out<=166;
				end
				if(in == 794) begin
					state<=3;
					out<=167;
				end
				if(in == 795) begin
					state<=3;
					out<=168;
				end
				if(in == 796) begin
					state<=3;
					out<=169;
				end
				if(in == 797) begin
					state<=3;
					out<=170;
				end
				if(in == 798) begin
					state<=3;
					out<=171;
				end
				if(in == 799) begin
					state<=3;
					out<=172;
				end
				if(in == 800) begin
					state<=3;
					out<=173;
				end
				if(in == 801) begin
					state<=14;
					out<=174;
				end
				if(in == 802) begin
					state<=14;
					out<=175;
				end
				if(in == 803) begin
					state<=14;
					out<=176;
				end
				if(in == 804) begin
					state<=14;
					out<=177;
				end
				if(in == 805) begin
					state<=14;
					out<=178;
				end
				if(in == 806) begin
					state<=14;
					out<=179;
				end
				if(in == 807) begin
					state<=3;
					out<=180;
				end
				if(in == 808) begin
					state<=3;
					out<=181;
				end
				if(in == 809) begin
					state<=3;
					out<=182;
				end
				if(in == 810) begin
					state<=3;
					out<=183;
				end
				if(in == 811) begin
					state<=3;
					out<=184;
				end
				if(in == 812) begin
					state<=3;
					out<=185;
				end
				if(in == 813) begin
					state<=14;
					out<=186;
				end
				if(in == 814) begin
					state<=14;
					out<=187;
				end
				if(in == 815) begin
					state<=14;
					out<=188;
				end
				if(in == 816) begin
					state<=14;
					out<=189;
				end
				if(in == 817) begin
					state<=14;
					out<=190;
				end
				if(in == 818) begin
					state<=14;
					out<=191;
				end
				if(in == 819) begin
					state<=14;
					out<=192;
				end
				if(in == 820) begin
					state<=14;
					out<=193;
				end
				if(in == 821) begin
					state<=14;
					out<=194;
				end
				if(in == 822) begin
					state<=14;
					out<=195;
				end
				if(in == 823) begin
					state<=14;
					out<=196;
				end
				if(in == 824) begin
					state<=14;
					out<=197;
				end
				if(in == 825) begin
					state<=14;
					out<=198;
				end
				if(in == 826) begin
					state<=14;
					out<=199;
				end
				if(in == 827) begin
					state<=14;
					out<=200;
				end
				if(in == 828) begin
					state<=14;
					out<=201;
				end
				if(in == 829) begin
					state<=14;
					out<=202;
				end
				if(in == 830) begin
					state<=14;
					out<=203;
				end
				if(in == 831) begin
					state<=14;
					out<=204;
				end
				if(in == 832) begin
					state<=14;
					out<=205;
				end
				if(in == 833) begin
					state<=14;
					out<=206;
				end
				if(in == 834) begin
					state<=14;
					out<=207;
				end
				if(in == 835) begin
					state<=14;
					out<=208;
				end
				if(in == 836) begin
					state<=14;
					out<=209;
				end
				if(in == 837) begin
					state<=14;
					out<=210;
				end
				if(in == 838) begin
					state<=14;
					out<=211;
				end
				if(in == 839) begin
					state<=14;
					out<=212;
				end
				if(in == 840) begin
					state<=14;
					out<=213;
				end
				if(in == 841) begin
					state<=14;
					out<=214;
				end
				if(in == 842) begin
					state<=14;
					out<=215;
				end
				if(in == 843) begin
					state<=14;
					out<=216;
				end
				if(in == 844) begin
					state<=14;
					out<=217;
				end
				if(in == 845) begin
					state<=14;
					out<=218;
				end
				if(in == 846) begin
					state<=14;
					out<=219;
				end
				if(in == 847) begin
					state<=14;
					out<=220;
				end
				if(in == 848) begin
					state<=14;
					out<=221;
				end
				if(in == 849) begin
					state<=14;
					out<=222;
				end
				if(in == 850) begin
					state<=14;
					out<=223;
				end
				if(in == 851) begin
					state<=14;
					out<=224;
				end
				if(in == 852) begin
					state<=14;
					out<=225;
				end
				if(in == 853) begin
					state<=14;
					out<=226;
				end
				if(in == 854) begin
					state<=14;
					out<=227;
				end
				if(in == 855) begin
					state<=14;
					out<=228;
				end
				if(in == 856) begin
					state<=14;
					out<=229;
				end
				if(in == 857) begin
					state<=14;
					out<=230;
				end
				if(in == 858) begin
					state<=14;
					out<=231;
				end
				if(in == 859) begin
					state<=14;
					out<=232;
				end
				if(in == 860) begin
					state<=14;
					out<=233;
				end
				if(in == 861) begin
					state<=14;
					out<=234;
				end
				if(in == 862) begin
					state<=14;
					out<=235;
				end
				if(in == 863) begin
					state<=14;
					out<=236;
				end
				if(in == 864) begin
					state<=14;
					out<=237;
				end
				if(in == 865) begin
					state<=3;
					out<=238;
				end
				if(in == 866) begin
					state<=3;
					out<=239;
				end
				if(in == 867) begin
					state<=3;
					out<=240;
				end
				if(in == 868) begin
					state<=3;
					out<=241;
				end
				if(in == 869) begin
					state<=3;
					out<=242;
				end
				if(in == 870) begin
					state<=3;
					out<=243;
				end
				if(in == 871) begin
					state<=3;
					out<=244;
				end
				if(in == 872) begin
					state<=3;
					out<=245;
				end
				if(in == 873) begin
					state<=3;
					out<=246;
				end
				if(in == 874) begin
					state<=3;
					out<=247;
				end
				if(in == 875) begin
					state<=3;
					out<=248;
				end
				if(in == 876) begin
					state<=3;
					out<=249;
				end
				if(in == 877) begin
					state<=3;
					out<=250;
				end
				if(in == 878) begin
					state<=3;
					out<=251;
				end
				if(in == 879) begin
					state<=3;
					out<=252;
				end
				if(in == 880) begin
					state<=3;
					out<=253;
				end
				if(in == 881) begin
					state<=3;
					out<=254;
				end
				if(in == 882) begin
					state<=3;
					out<=255;
				end
				if(in == 883) begin
					state<=3;
					out<=0;
				end
				if(in == 884) begin
					state<=3;
					out<=1;
				end
				if(in == 885) begin
					state<=3;
					out<=2;
				end
				if(in == 886) begin
					state<=3;
					out<=3;
				end
				if(in == 887) begin
					state<=3;
					out<=4;
				end
				if(in == 888) begin
					state<=3;
					out<=5;
				end
				if(in == 889) begin
					state<=3;
					out<=6;
				end
				if(in == 890) begin
					state<=3;
					out<=7;
				end
				if(in == 891) begin
					state<=3;
					out<=8;
				end
				if(in == 892) begin
					state<=3;
					out<=9;
				end
				if(in == 893) begin
					state<=3;
					out<=10;
				end
				if(in == 894) begin
					state<=3;
					out<=11;
				end
				if(in == 895) begin
					state<=3;
					out<=12;
				end
				if(in == 896) begin
					state<=3;
					out<=13;
				end
				if(in == 897) begin
					state<=3;
					out<=14;
				end
				if(in == 898) begin
					state<=3;
					out<=15;
				end
				if(in == 899) begin
					state<=3;
					out<=16;
				end
				if(in == 900) begin
					state<=3;
					out<=17;
				end
				if(in == 901) begin
					state<=3;
					out<=18;
				end
				if(in == 902) begin
					state<=3;
					out<=19;
				end
				if(in == 903) begin
					state<=3;
					out<=20;
				end
				if(in == 904) begin
					state<=3;
					out<=21;
				end
				if(in == 905) begin
					state<=3;
					out<=22;
				end
				if(in == 906) begin
					state<=3;
					out<=23;
				end
				if(in == 907) begin
					state<=3;
					out<=24;
				end
				if(in == 908) begin
					state<=3;
					out<=25;
				end
				if(in == 909) begin
					state<=3;
					out<=26;
				end
				if(in == 910) begin
					state<=3;
					out<=27;
				end
				if(in == 911) begin
					state<=3;
					out<=28;
				end
				if(in == 912) begin
					state<=3;
					out<=29;
				end
				if(in == 913) begin
					state<=3;
					out<=30;
				end
				if(in == 914) begin
					state<=3;
					out<=31;
				end
				if(in == 915) begin
					state<=3;
					out<=32;
				end
				if(in == 916) begin
					state<=3;
					out<=33;
				end
				if(in == 917) begin
					state<=14;
					out<=34;
				end
				if(in == 918) begin
					state<=14;
					out<=35;
				end
				if(in == 919) begin
					state<=14;
					out<=36;
				end
				if(in == 920) begin
					state<=14;
					out<=37;
				end
				if(in == 921) begin
					state<=14;
					out<=38;
				end
				if(in == 922) begin
					state<=14;
					out<=39;
				end
				if(in == 923) begin
					state<=3;
					out<=40;
				end
				if(in == 924) begin
					state<=3;
					out<=41;
				end
				if(in == 925) begin
					state<=3;
					out<=42;
				end
				if(in == 926) begin
					state<=3;
					out<=43;
				end
				if(in == 927) begin
					state<=3;
					out<=44;
				end
				if(in == 928) begin
					state<=3;
					out<=45;
				end
			end
			14: begin
				if(in == 0) begin
					state<=14;
					out<=46;
				end
				if(in == 1) begin
					state<=1;
					out<=47;
				end
				if(in == 2) begin
					state<=14;
					out<=48;
				end
				if(in == 3) begin
					state<=14;
					out<=49;
				end
				if(in == 4) begin
					state<=14;
					out<=50;
				end
				if(in == 5) begin
					state<=14;
					out<=51;
				end
				if(in == 6) begin
					state<=14;
					out<=52;
				end
				if(in == 7) begin
					state<=14;
					out<=53;
				end
				if(in == 8) begin
					state<=14;
					out<=54;
				end
				if(in == 9) begin
					state<=14;
					out<=55;
				end
				if(in == 10) begin
					state<=14;
					out<=56;
				end
				if(in == 11) begin
					state<=14;
					out<=57;
				end
				if(in == 12) begin
					state<=14;
					out<=58;
				end
				if(in == 13) begin
					state<=14;
					out<=59;
				end
				if(in == 14) begin
					state<=14;
					out<=60;
				end
				if(in == 15) begin
					state<=14;
					out<=61;
				end
				if(in == 16) begin
					state<=14;
					out<=62;
				end
				if(in == 17) begin
					state<=14;
					out<=63;
				end
				if(in == 18) begin
					state<=14;
					out<=64;
				end
				if(in == 19) begin
					state<=14;
					out<=65;
				end
				if(in == 20) begin
					state<=14;
					out<=66;
				end
				if(in == 21) begin
					state<=14;
					out<=67;
				end
				if(in == 22) begin
					state<=14;
					out<=68;
				end
				if(in == 23) begin
					state<=14;
					out<=69;
				end
				if(in == 24) begin
					state<=14;
					out<=70;
				end
				if(in == 25) begin
					state<=14;
					out<=71;
				end
				if(in == 26) begin
					state<=14;
					out<=72;
				end
				if(in == 27) begin
					state<=14;
					out<=73;
				end
				if(in == 28) begin
					state<=14;
					out<=74;
				end
				if(in == 29) begin
					state<=14;
					out<=75;
				end
				if(in == 30) begin
					state<=14;
					out<=76;
				end
				if(in == 31) begin
					state<=14;
					out<=77;
				end
				if(in == 32) begin
					state<=14;
					out<=78;
				end
				if(in == 33) begin
					state<=14;
					out<=79;
				end
				if(in == 34) begin
					state<=14;
					out<=80;
				end
				if(in == 35) begin
					state<=14;
					out<=81;
				end
				if(in == 36) begin
					state<=14;
					out<=82;
				end
				if(in == 37) begin
					state<=14;
					out<=83;
				end
				if(in == 38) begin
					state<=14;
					out<=84;
				end
				if(in == 39) begin
					state<=14;
					out<=85;
				end
				if(in == 40) begin
					state<=14;
					out<=86;
				end
				if(in == 41) begin
					state<=14;
					out<=87;
				end
				if(in == 42) begin
					state<=14;
					out<=88;
				end
				if(in == 43) begin
					state<=14;
					out<=89;
				end
				if(in == 44) begin
					state<=14;
					out<=90;
				end
				if(in == 45) begin
					state<=14;
					out<=91;
				end
				if(in == 46) begin
					state<=14;
					out<=92;
				end
				if(in == 47) begin
					state<=14;
					out<=93;
				end
				if(in == 48) begin
					state<=14;
					out<=94;
				end
				if(in == 49) begin
					state<=14;
					out<=95;
				end
				if(in == 50) begin
					state<=14;
					out<=96;
				end
				if(in == 51) begin
					state<=14;
					out<=97;
				end
				if(in == 52) begin
					state<=14;
					out<=98;
				end
				if(in == 53) begin
					state<=14;
					out<=99;
				end
				if(in == 54) begin
					state<=14;
					out<=100;
				end
				if(in == 55) begin
					state<=14;
					out<=101;
				end
				if(in == 56) begin
					state<=14;
					out<=102;
				end
				if(in == 57) begin
					state<=14;
					out<=103;
				end
				if(in == 58) begin
					state<=14;
					out<=104;
				end
				if(in == 59) begin
					state<=14;
					out<=105;
				end
				if(in == 60) begin
					state<=14;
					out<=106;
				end
				if(in == 61) begin
					state<=14;
					out<=107;
				end
				if(in == 62) begin
					state<=14;
					out<=108;
				end
				if(in == 63) begin
					state<=14;
					out<=109;
				end
				if(in == 64) begin
					state<=14;
					out<=110;
				end
				if(in == 65) begin
					state<=14;
					out<=111;
				end
				if(in == 66) begin
					state<=14;
					out<=112;
				end
				if(in == 67) begin
					state<=14;
					out<=113;
				end
				if(in == 68) begin
					state<=14;
					out<=114;
				end
				if(in == 69) begin
					state<=14;
					out<=115;
				end
				if(in == 70) begin
					state<=14;
					out<=116;
				end
				if(in == 71) begin
					state<=14;
					out<=117;
				end
				if(in == 72) begin
					state<=14;
					out<=118;
				end
				if(in == 73) begin
					state<=14;
					out<=119;
				end
				if(in == 74) begin
					state<=14;
					out<=120;
				end
				if(in == 75) begin
					state<=14;
					out<=121;
				end
				if(in == 76) begin
					state<=14;
					out<=122;
				end
				if(in == 77) begin
					state<=14;
					out<=123;
				end
				if(in == 78) begin
					state<=14;
					out<=124;
				end
				if(in == 79) begin
					state<=14;
					out<=125;
				end
				if(in == 80) begin
					state<=14;
					out<=126;
				end
				if(in == 81) begin
					state<=14;
					out<=127;
				end
				if(in == 82) begin
					state<=14;
					out<=128;
				end
				if(in == 83) begin
					state<=14;
					out<=129;
				end
				if(in == 84) begin
					state<=14;
					out<=130;
				end
				if(in == 85) begin
					state<=14;
					out<=131;
				end
				if(in == 86) begin
					state<=14;
					out<=132;
				end
				if(in == 87) begin
					state<=14;
					out<=133;
				end
				if(in == 88) begin
					state<=14;
					out<=134;
				end
				if(in == 89) begin
					state<=14;
					out<=135;
				end
				if(in == 90) begin
					state<=14;
					out<=136;
				end
				if(in == 91) begin
					state<=14;
					out<=137;
				end
				if(in == 92) begin
					state<=14;
					out<=138;
				end
				if(in == 93) begin
					state<=14;
					out<=139;
				end
				if(in == 94) begin
					state<=14;
					out<=140;
				end
				if(in == 95) begin
					state<=14;
					out<=141;
				end
				if(in == 96) begin
					state<=14;
					out<=142;
				end
				if(in == 97) begin
					state<=14;
					out<=143;
				end
				if(in == 98) begin
					state<=14;
					out<=144;
				end
				if(in == 99) begin
					state<=14;
					out<=145;
				end
				if(in == 100) begin
					state<=14;
					out<=146;
				end
				if(in == 101) begin
					state<=14;
					out<=147;
				end
				if(in == 102) begin
					state<=14;
					out<=148;
				end
				if(in == 103) begin
					state<=14;
					out<=149;
				end
				if(in == 104) begin
					state<=14;
					out<=150;
				end
				if(in == 105) begin
					state<=14;
					out<=151;
				end
				if(in == 106) begin
					state<=14;
					out<=152;
				end
				if(in == 107) begin
					state<=14;
					out<=153;
				end
				if(in == 108) begin
					state<=14;
					out<=154;
				end
				if(in == 109) begin
					state<=14;
					out<=155;
				end
				if(in == 110) begin
					state<=14;
					out<=156;
				end
				if(in == 111) begin
					state<=14;
					out<=157;
				end
				if(in == 112) begin
					state<=14;
					out<=158;
				end
				if(in == 113) begin
					state<=14;
					out<=159;
				end
				if(in == 114) begin
					state<=14;
					out<=160;
				end
				if(in == 115) begin
					state<=14;
					out<=161;
				end
				if(in == 116) begin
					state<=14;
					out<=162;
				end
				if(in == 117) begin
					state<=1;
					out<=163;
				end
				if(in == 118) begin
					state<=1;
					out<=164;
				end
				if(in == 119) begin
					state<=1;
					out<=165;
				end
				if(in == 120) begin
					state<=1;
					out<=166;
				end
				if(in == 121) begin
					state<=1;
					out<=167;
				end
				if(in == 122) begin
					state<=1;
					out<=168;
				end
				if(in == 123) begin
					state<=1;
					out<=169;
				end
				if(in == 124) begin
					state<=1;
					out<=170;
				end
				if(in == 125) begin
					state<=1;
					out<=171;
				end
				if(in == 126) begin
					state<=1;
					out<=172;
				end
				if(in == 127) begin
					state<=1;
					out<=173;
				end
				if(in == 128) begin
					state<=1;
					out<=174;
				end
				if(in == 129) begin
					state<=1;
					out<=175;
				end
				if(in == 130) begin
					state<=1;
					out<=176;
				end
				if(in == 131) begin
					state<=1;
					out<=177;
				end
				if(in == 132) begin
					state<=1;
					out<=178;
				end
				if(in == 133) begin
					state<=1;
					out<=179;
				end
				if(in == 134) begin
					state<=1;
					out<=180;
				end
				if(in == 135) begin
					state<=1;
					out<=181;
				end
				if(in == 136) begin
					state<=1;
					out<=182;
				end
				if(in == 137) begin
					state<=1;
					out<=183;
				end
				if(in == 138) begin
					state<=1;
					out<=184;
				end
				if(in == 139) begin
					state<=1;
					out<=185;
				end
				if(in == 140) begin
					state<=1;
					out<=186;
				end
				if(in == 141) begin
					state<=1;
					out<=187;
				end
				if(in == 142) begin
					state<=1;
					out<=188;
				end
				if(in == 143) begin
					state<=1;
					out<=189;
				end
				if(in == 144) begin
					state<=1;
					out<=190;
				end
				if(in == 145) begin
					state<=1;
					out<=191;
				end
				if(in == 146) begin
					state<=1;
					out<=192;
				end
				if(in == 147) begin
					state<=1;
					out<=193;
				end
				if(in == 148) begin
					state<=1;
					out<=194;
				end
				if(in == 149) begin
					state<=1;
					out<=195;
				end
				if(in == 150) begin
					state<=1;
					out<=196;
				end
				if(in == 151) begin
					state<=1;
					out<=197;
				end
				if(in == 152) begin
					state<=1;
					out<=198;
				end
				if(in == 153) begin
					state<=1;
					out<=199;
				end
				if(in == 154) begin
					state<=1;
					out<=200;
				end
				if(in == 155) begin
					state<=1;
					out<=201;
				end
				if(in == 156) begin
					state<=1;
					out<=202;
				end
				if(in == 157) begin
					state<=1;
					out<=203;
				end
				if(in == 158) begin
					state<=1;
					out<=204;
				end
				if(in == 159) begin
					state<=1;
					out<=205;
				end
				if(in == 160) begin
					state<=1;
					out<=206;
				end
				if(in == 161) begin
					state<=1;
					out<=207;
				end
				if(in == 162) begin
					state<=1;
					out<=208;
				end
				if(in == 163) begin
					state<=1;
					out<=209;
				end
				if(in == 164) begin
					state<=1;
					out<=210;
				end
				if(in == 165) begin
					state<=1;
					out<=211;
				end
				if(in == 166) begin
					state<=1;
					out<=212;
				end
				if(in == 167) begin
					state<=1;
					out<=213;
				end
				if(in == 168) begin
					state<=1;
					out<=214;
				end
				if(in == 169) begin
					state<=1;
					out<=215;
				end
				if(in == 170) begin
					state<=1;
					out<=216;
				end
				if(in == 171) begin
					state<=1;
					out<=217;
				end
				if(in == 172) begin
					state<=1;
					out<=218;
				end
				if(in == 173) begin
					state<=1;
					out<=219;
				end
				if(in == 174) begin
					state<=1;
					out<=220;
				end
				if(in == 175) begin
					state<=1;
					out<=221;
				end
				if(in == 176) begin
					state<=1;
					out<=222;
				end
				if(in == 177) begin
					state<=1;
					out<=223;
				end
				if(in == 178) begin
					state<=1;
					out<=224;
				end
				if(in == 179) begin
					state<=1;
					out<=225;
				end
				if(in == 180) begin
					state<=1;
					out<=226;
				end
				if(in == 181) begin
					state<=1;
					out<=227;
				end
				if(in == 182) begin
					state<=1;
					out<=228;
				end
				if(in == 183) begin
					state<=1;
					out<=229;
				end
				if(in == 184) begin
					state<=1;
					out<=230;
				end
				if(in == 185) begin
					state<=1;
					out<=231;
				end
				if(in == 186) begin
					state<=1;
					out<=232;
				end
				if(in == 187) begin
					state<=1;
					out<=233;
				end
				if(in == 188) begin
					state<=1;
					out<=234;
				end
				if(in == 189) begin
					state<=1;
					out<=235;
				end
				if(in == 190) begin
					state<=1;
					out<=236;
				end
				if(in == 191) begin
					state<=1;
					out<=237;
				end
				if(in == 192) begin
					state<=1;
					out<=238;
				end
				if(in == 193) begin
					state<=1;
					out<=239;
				end
				if(in == 194) begin
					state<=1;
					out<=240;
				end
				if(in == 195) begin
					state<=1;
					out<=241;
				end
				if(in == 196) begin
					state<=1;
					out<=242;
				end
				if(in == 197) begin
					state<=1;
					out<=243;
				end
				if(in == 198) begin
					state<=1;
					out<=244;
				end
				if(in == 199) begin
					state<=1;
					out<=245;
				end
				if(in == 200) begin
					state<=1;
					out<=246;
				end
				if(in == 201) begin
					state<=1;
					out<=247;
				end
				if(in == 202) begin
					state<=1;
					out<=248;
				end
				if(in == 203) begin
					state<=1;
					out<=249;
				end
				if(in == 204) begin
					state<=1;
					out<=250;
				end
				if(in == 205) begin
					state<=1;
					out<=251;
				end
				if(in == 206) begin
					state<=1;
					out<=252;
				end
				if(in == 207) begin
					state<=1;
					out<=253;
				end
				if(in == 208) begin
					state<=1;
					out<=254;
				end
				if(in == 209) begin
					state<=1;
					out<=255;
				end
				if(in == 210) begin
					state<=1;
					out<=0;
				end
				if(in == 211) begin
					state<=1;
					out<=1;
				end
				if(in == 212) begin
					state<=1;
					out<=2;
				end
				if(in == 213) begin
					state<=1;
					out<=3;
				end
				if(in == 214) begin
					state<=1;
					out<=4;
				end
				if(in == 215) begin
					state<=1;
					out<=5;
				end
				if(in == 216) begin
					state<=1;
					out<=6;
				end
				if(in == 217) begin
					state<=1;
					out<=7;
				end
				if(in == 218) begin
					state<=1;
					out<=8;
				end
				if(in == 219) begin
					state<=1;
					out<=9;
				end
				if(in == 220) begin
					state<=1;
					out<=10;
				end
				if(in == 221) begin
					state<=1;
					out<=11;
				end
				if(in == 222) begin
					state<=1;
					out<=12;
				end
				if(in == 223) begin
					state<=1;
					out<=13;
				end
				if(in == 224) begin
					state<=1;
					out<=14;
				end
				if(in == 225) begin
					state<=1;
					out<=15;
				end
				if(in == 226) begin
					state<=1;
					out<=16;
				end
				if(in == 227) begin
					state<=1;
					out<=17;
				end
				if(in == 228) begin
					state<=1;
					out<=18;
				end
				if(in == 229) begin
					state<=1;
					out<=19;
				end
				if(in == 230) begin
					state<=1;
					out<=20;
				end
				if(in == 231) begin
					state<=1;
					out<=21;
				end
				if(in == 232) begin
					state<=1;
					out<=22;
				end
				if(in == 233) begin
					state<=15;
					out<=23;
				end
				if(in == 234) begin
					state<=15;
					out<=24;
				end
				if(in == 235) begin
					state<=15;
					out<=25;
				end
				if(in == 236) begin
					state<=15;
					out<=26;
				end
				if(in == 237) begin
					state<=15;
					out<=27;
				end
				if(in == 238) begin
					state<=15;
					out<=28;
				end
				if(in == 239) begin
					state<=15;
					out<=29;
				end
				if(in == 240) begin
					state<=15;
					out<=30;
				end
				if(in == 241) begin
					state<=15;
					out<=31;
				end
				if(in == 242) begin
					state<=15;
					out<=32;
				end
				if(in == 243) begin
					state<=15;
					out<=33;
				end
				if(in == 244) begin
					state<=15;
					out<=34;
				end
				if(in == 245) begin
					state<=15;
					out<=35;
				end
				if(in == 246) begin
					state<=15;
					out<=36;
				end
				if(in == 247) begin
					state<=15;
					out<=37;
				end
				if(in == 248) begin
					state<=15;
					out<=38;
				end
				if(in == 249) begin
					state<=15;
					out<=39;
				end
				if(in == 250) begin
					state<=15;
					out<=40;
				end
				if(in == 251) begin
					state<=15;
					out<=41;
				end
				if(in == 252) begin
					state<=15;
					out<=42;
				end
				if(in == 253) begin
					state<=15;
					out<=43;
				end
				if(in == 254) begin
					state<=15;
					out<=44;
				end
				if(in == 255) begin
					state<=15;
					out<=45;
				end
				if(in == 256) begin
					state<=15;
					out<=46;
				end
				if(in == 257) begin
					state<=15;
					out<=47;
				end
				if(in == 258) begin
					state<=15;
					out<=48;
				end
				if(in == 259) begin
					state<=15;
					out<=49;
				end
				if(in == 260) begin
					state<=15;
					out<=50;
				end
				if(in == 261) begin
					state<=15;
					out<=51;
				end
				if(in == 262) begin
					state<=15;
					out<=52;
				end
				if(in == 263) begin
					state<=15;
					out<=53;
				end
				if(in == 264) begin
					state<=15;
					out<=54;
				end
				if(in == 265) begin
					state<=15;
					out<=55;
				end
				if(in == 266) begin
					state<=15;
					out<=56;
				end
				if(in == 267) begin
					state<=15;
					out<=57;
				end
				if(in == 268) begin
					state<=15;
					out<=58;
				end
				if(in == 269) begin
					state<=15;
					out<=59;
				end
				if(in == 270) begin
					state<=15;
					out<=60;
				end
				if(in == 271) begin
					state<=15;
					out<=61;
				end
				if(in == 272) begin
					state<=15;
					out<=62;
				end
				if(in == 273) begin
					state<=15;
					out<=63;
				end
				if(in == 274) begin
					state<=15;
					out<=64;
				end
				if(in == 275) begin
					state<=15;
					out<=65;
				end
				if(in == 276) begin
					state<=15;
					out<=66;
				end
				if(in == 277) begin
					state<=15;
					out<=67;
				end
				if(in == 278) begin
					state<=15;
					out<=68;
				end
				if(in == 279) begin
					state<=15;
					out<=69;
				end
				if(in == 280) begin
					state<=15;
					out<=70;
				end
				if(in == 281) begin
					state<=15;
					out<=71;
				end
				if(in == 282) begin
					state<=15;
					out<=72;
				end
				if(in == 283) begin
					state<=15;
					out<=73;
				end
				if(in == 284) begin
					state<=15;
					out<=74;
				end
				if(in == 285) begin
					state<=15;
					out<=75;
				end
				if(in == 286) begin
					state<=15;
					out<=76;
				end
				if(in == 287) begin
					state<=15;
					out<=77;
				end
				if(in == 288) begin
					state<=15;
					out<=78;
				end
				if(in == 289) begin
					state<=15;
					out<=79;
				end
				if(in == 290) begin
					state<=15;
					out<=80;
				end
				if(in == 291) begin
					state<=15;
					out<=81;
				end
				if(in == 292) begin
					state<=15;
					out<=82;
				end
				if(in == 293) begin
					state<=15;
					out<=83;
				end
				if(in == 294) begin
					state<=15;
					out<=84;
				end
				if(in == 295) begin
					state<=15;
					out<=85;
				end
				if(in == 296) begin
					state<=15;
					out<=86;
				end
				if(in == 297) begin
					state<=15;
					out<=87;
				end
				if(in == 298) begin
					state<=15;
					out<=88;
				end
				if(in == 299) begin
					state<=15;
					out<=89;
				end
				if(in == 300) begin
					state<=15;
					out<=90;
				end
				if(in == 301) begin
					state<=15;
					out<=91;
				end
				if(in == 302) begin
					state<=15;
					out<=92;
				end
				if(in == 303) begin
					state<=15;
					out<=93;
				end
				if(in == 304) begin
					state<=15;
					out<=94;
				end
				if(in == 305) begin
					state<=15;
					out<=95;
				end
				if(in == 306) begin
					state<=15;
					out<=96;
				end
				if(in == 307) begin
					state<=15;
					out<=97;
				end
				if(in == 308) begin
					state<=15;
					out<=98;
				end
				if(in == 309) begin
					state<=15;
					out<=99;
				end
				if(in == 310) begin
					state<=15;
					out<=100;
				end
				if(in == 311) begin
					state<=15;
					out<=101;
				end
				if(in == 312) begin
					state<=15;
					out<=102;
				end
				if(in == 313) begin
					state<=15;
					out<=103;
				end
				if(in == 314) begin
					state<=15;
					out<=104;
				end
				if(in == 315) begin
					state<=15;
					out<=105;
				end
				if(in == 316) begin
					state<=15;
					out<=106;
				end
				if(in == 317) begin
					state<=15;
					out<=107;
				end
				if(in == 318) begin
					state<=15;
					out<=108;
				end
				if(in == 319) begin
					state<=15;
					out<=109;
				end
				if(in == 320) begin
					state<=15;
					out<=110;
				end
				if(in == 321) begin
					state<=15;
					out<=111;
				end
				if(in == 322) begin
					state<=15;
					out<=112;
				end
				if(in == 323) begin
					state<=15;
					out<=113;
				end
				if(in == 324) begin
					state<=15;
					out<=114;
				end
				if(in == 325) begin
					state<=15;
					out<=115;
				end
				if(in == 326) begin
					state<=15;
					out<=116;
				end
				if(in == 327) begin
					state<=15;
					out<=117;
				end
				if(in == 328) begin
					state<=15;
					out<=118;
				end
				if(in == 329) begin
					state<=15;
					out<=119;
				end
				if(in == 330) begin
					state<=15;
					out<=120;
				end
				if(in == 331) begin
					state<=15;
					out<=121;
				end
				if(in == 332) begin
					state<=15;
					out<=122;
				end
				if(in == 333) begin
					state<=15;
					out<=123;
				end
				if(in == 334) begin
					state<=15;
					out<=124;
				end
				if(in == 335) begin
					state<=15;
					out<=125;
				end
				if(in == 336) begin
					state<=15;
					out<=126;
				end
				if(in == 337) begin
					state<=15;
					out<=127;
				end
				if(in == 338) begin
					state<=15;
					out<=128;
				end
				if(in == 339) begin
					state<=15;
					out<=129;
				end
				if(in == 340) begin
					state<=15;
					out<=130;
				end
				if(in == 341) begin
					state<=15;
					out<=131;
				end
				if(in == 342) begin
					state<=15;
					out<=132;
				end
				if(in == 343) begin
					state<=15;
					out<=133;
				end
				if(in == 344) begin
					state<=15;
					out<=134;
				end
				if(in == 345) begin
					state<=15;
					out<=135;
				end
				if(in == 346) begin
					state<=15;
					out<=136;
				end
				if(in == 347) begin
					state<=15;
					out<=137;
				end
				if(in == 348) begin
					state<=15;
					out<=138;
				end
				if(in == 349) begin
					state<=16;
					out<=139;
				end
				if(in == 350) begin
					state<=16;
					out<=140;
				end
				if(in == 351) begin
					state<=16;
					out<=141;
				end
				if(in == 352) begin
					state<=16;
					out<=142;
				end
				if(in == 353) begin
					state<=16;
					out<=143;
				end
				if(in == 354) begin
					state<=16;
					out<=144;
				end
				if(in == 355) begin
					state<=16;
					out<=145;
				end
				if(in == 356) begin
					state<=16;
					out<=146;
				end
				if(in == 357) begin
					state<=16;
					out<=147;
				end
				if(in == 358) begin
					state<=16;
					out<=148;
				end
				if(in == 359) begin
					state<=16;
					out<=149;
				end
				if(in == 360) begin
					state<=16;
					out<=150;
				end
				if(in == 361) begin
					state<=16;
					out<=151;
				end
				if(in == 362) begin
					state<=16;
					out<=152;
				end
				if(in == 363) begin
					state<=16;
					out<=153;
				end
				if(in == 364) begin
					state<=16;
					out<=154;
				end
				if(in == 365) begin
					state<=16;
					out<=155;
				end
				if(in == 366) begin
					state<=16;
					out<=156;
				end
				if(in == 367) begin
					state<=16;
					out<=157;
				end
				if(in == 368) begin
					state<=16;
					out<=158;
				end
				if(in == 369) begin
					state<=16;
					out<=159;
				end
				if(in == 370) begin
					state<=16;
					out<=160;
				end
				if(in == 371) begin
					state<=16;
					out<=161;
				end
				if(in == 372) begin
					state<=16;
					out<=162;
				end
				if(in == 373) begin
					state<=16;
					out<=163;
				end
				if(in == 374) begin
					state<=16;
					out<=164;
				end
				if(in == 375) begin
					state<=16;
					out<=165;
				end
				if(in == 376) begin
					state<=16;
					out<=166;
				end
				if(in == 377) begin
					state<=16;
					out<=167;
				end
				if(in == 378) begin
					state<=16;
					out<=168;
				end
				if(in == 379) begin
					state<=16;
					out<=169;
				end
				if(in == 380) begin
					state<=16;
					out<=170;
				end
				if(in == 381) begin
					state<=16;
					out<=171;
				end
				if(in == 382) begin
					state<=16;
					out<=172;
				end
				if(in == 383) begin
					state<=16;
					out<=173;
				end
				if(in == 384) begin
					state<=16;
					out<=174;
				end
				if(in == 385) begin
					state<=16;
					out<=175;
				end
				if(in == 386) begin
					state<=16;
					out<=176;
				end
				if(in == 387) begin
					state<=16;
					out<=177;
				end
				if(in == 388) begin
					state<=16;
					out<=178;
				end
				if(in == 389) begin
					state<=16;
					out<=179;
				end
				if(in == 390) begin
					state<=16;
					out<=180;
				end
				if(in == 391) begin
					state<=16;
					out<=181;
				end
				if(in == 392) begin
					state<=16;
					out<=182;
				end
				if(in == 393) begin
					state<=16;
					out<=183;
				end
				if(in == 394) begin
					state<=16;
					out<=184;
				end
				if(in == 395) begin
					state<=16;
					out<=185;
				end
				if(in == 396) begin
					state<=16;
					out<=186;
				end
				if(in == 397) begin
					state<=16;
					out<=187;
				end
				if(in == 398) begin
					state<=16;
					out<=188;
				end
				if(in == 399) begin
					state<=16;
					out<=189;
				end
				if(in == 400) begin
					state<=16;
					out<=190;
				end
				if(in == 401) begin
					state<=16;
					out<=191;
				end
				if(in == 402) begin
					state<=16;
					out<=192;
				end
				if(in == 403) begin
					state<=16;
					out<=193;
				end
				if(in == 404) begin
					state<=16;
					out<=194;
				end
				if(in == 405) begin
					state<=16;
					out<=195;
				end
				if(in == 406) begin
					state<=16;
					out<=196;
				end
				if(in == 407) begin
					state<=16;
					out<=197;
				end
				if(in == 408) begin
					state<=16;
					out<=198;
				end
				if(in == 409) begin
					state<=16;
					out<=199;
				end
				if(in == 410) begin
					state<=16;
					out<=200;
				end
				if(in == 411) begin
					state<=16;
					out<=201;
				end
				if(in == 412) begin
					state<=16;
					out<=202;
				end
				if(in == 413) begin
					state<=16;
					out<=203;
				end
				if(in == 414) begin
					state<=16;
					out<=204;
				end
				if(in == 415) begin
					state<=16;
					out<=205;
				end
				if(in == 416) begin
					state<=16;
					out<=206;
				end
				if(in == 417) begin
					state<=16;
					out<=207;
				end
				if(in == 418) begin
					state<=16;
					out<=208;
				end
				if(in == 419) begin
					state<=16;
					out<=209;
				end
				if(in == 420) begin
					state<=16;
					out<=210;
				end
				if(in == 421) begin
					state<=16;
					out<=211;
				end
				if(in == 422) begin
					state<=16;
					out<=212;
				end
				if(in == 423) begin
					state<=16;
					out<=213;
				end
				if(in == 424) begin
					state<=16;
					out<=214;
				end
				if(in == 425) begin
					state<=16;
					out<=215;
				end
				if(in == 426) begin
					state<=16;
					out<=216;
				end
				if(in == 427) begin
					state<=16;
					out<=217;
				end
				if(in == 428) begin
					state<=16;
					out<=218;
				end
				if(in == 429) begin
					state<=16;
					out<=219;
				end
				if(in == 430) begin
					state<=16;
					out<=220;
				end
				if(in == 431) begin
					state<=16;
					out<=221;
				end
				if(in == 432) begin
					state<=16;
					out<=222;
				end
				if(in == 433) begin
					state<=16;
					out<=223;
				end
				if(in == 434) begin
					state<=16;
					out<=224;
				end
				if(in == 435) begin
					state<=16;
					out<=225;
				end
				if(in == 436) begin
					state<=16;
					out<=226;
				end
				if(in == 437) begin
					state<=16;
					out<=227;
				end
				if(in == 438) begin
					state<=16;
					out<=228;
				end
				if(in == 439) begin
					state<=16;
					out<=229;
				end
				if(in == 440) begin
					state<=16;
					out<=230;
				end
				if(in == 441) begin
					state<=16;
					out<=231;
				end
				if(in == 442) begin
					state<=16;
					out<=232;
				end
				if(in == 443) begin
					state<=16;
					out<=233;
				end
				if(in == 444) begin
					state<=16;
					out<=234;
				end
				if(in == 445) begin
					state<=16;
					out<=235;
				end
				if(in == 446) begin
					state<=16;
					out<=236;
				end
				if(in == 447) begin
					state<=16;
					out<=237;
				end
				if(in == 448) begin
					state<=16;
					out<=238;
				end
				if(in == 449) begin
					state<=16;
					out<=239;
				end
				if(in == 450) begin
					state<=16;
					out<=240;
				end
				if(in == 451) begin
					state<=16;
					out<=241;
				end
				if(in == 452) begin
					state<=16;
					out<=242;
				end
				if(in == 453) begin
					state<=16;
					out<=243;
				end
				if(in == 454) begin
					state<=16;
					out<=244;
				end
				if(in == 455) begin
					state<=16;
					out<=245;
				end
				if(in == 456) begin
					state<=16;
					out<=246;
				end
				if(in == 457) begin
					state<=16;
					out<=247;
				end
				if(in == 458) begin
					state<=16;
					out<=248;
				end
				if(in == 459) begin
					state<=16;
					out<=249;
				end
				if(in == 460) begin
					state<=16;
					out<=250;
				end
				if(in == 461) begin
					state<=16;
					out<=251;
				end
				if(in == 462) begin
					state<=16;
					out<=252;
				end
				if(in == 463) begin
					state<=16;
					out<=253;
				end
				if(in == 464) begin
					state<=16;
					out<=254;
				end
				if(in == 465) begin
					state<=14;
					out<=255;
				end
				if(in == 466) begin
					state<=14;
					out<=0;
				end
				if(in == 467) begin
					state<=14;
					out<=1;
				end
				if(in == 468) begin
					state<=14;
					out<=2;
				end
				if(in == 469) begin
					state<=14;
					out<=3;
				end
				if(in == 470) begin
					state<=14;
					out<=4;
				end
				if(in == 471) begin
					state<=14;
					out<=5;
				end
				if(in == 472) begin
					state<=14;
					out<=6;
				end
				if(in == 473) begin
					state<=14;
					out<=7;
				end
				if(in == 474) begin
					state<=14;
					out<=8;
				end
				if(in == 475) begin
					state<=14;
					out<=9;
				end
				if(in == 476) begin
					state<=14;
					out<=10;
				end
				if(in == 477) begin
					state<=14;
					out<=11;
				end
				if(in == 478) begin
					state<=14;
					out<=12;
				end
				if(in == 479) begin
					state<=14;
					out<=13;
				end
				if(in == 480) begin
					state<=14;
					out<=14;
				end
				if(in == 481) begin
					state<=14;
					out<=15;
				end
				if(in == 482) begin
					state<=14;
					out<=16;
				end
				if(in == 483) begin
					state<=14;
					out<=17;
				end
				if(in == 484) begin
					state<=14;
					out<=18;
				end
				if(in == 485) begin
					state<=14;
					out<=19;
				end
				if(in == 486) begin
					state<=14;
					out<=20;
				end
				if(in == 487) begin
					state<=14;
					out<=21;
				end
				if(in == 488) begin
					state<=14;
					out<=22;
				end
				if(in == 489) begin
					state<=14;
					out<=23;
				end
				if(in == 490) begin
					state<=14;
					out<=24;
				end
				if(in == 491) begin
					state<=14;
					out<=25;
				end
				if(in == 492) begin
					state<=14;
					out<=26;
				end
				if(in == 493) begin
					state<=14;
					out<=27;
				end
				if(in == 494) begin
					state<=14;
					out<=28;
				end
				if(in == 495) begin
					state<=14;
					out<=29;
				end
				if(in == 496) begin
					state<=14;
					out<=30;
				end
				if(in == 497) begin
					state<=14;
					out<=31;
				end
				if(in == 498) begin
					state<=14;
					out<=32;
				end
				if(in == 499) begin
					state<=14;
					out<=33;
				end
				if(in == 500) begin
					state<=14;
					out<=34;
				end
				if(in == 501) begin
					state<=14;
					out<=35;
				end
				if(in == 502) begin
					state<=14;
					out<=36;
				end
				if(in == 503) begin
					state<=14;
					out<=37;
				end
				if(in == 504) begin
					state<=14;
					out<=38;
				end
				if(in == 505) begin
					state<=14;
					out<=39;
				end
				if(in == 506) begin
					state<=14;
					out<=40;
				end
				if(in == 507) begin
					state<=14;
					out<=41;
				end
				if(in == 508) begin
					state<=14;
					out<=42;
				end
				if(in == 509) begin
					state<=14;
					out<=43;
				end
				if(in == 510) begin
					state<=14;
					out<=44;
				end
				if(in == 511) begin
					state<=14;
					out<=45;
				end
				if(in == 512) begin
					state<=14;
					out<=46;
				end
				if(in == 513) begin
					state<=14;
					out<=47;
				end
				if(in == 514) begin
					state<=14;
					out<=48;
				end
				if(in == 515) begin
					state<=14;
					out<=49;
				end
				if(in == 516) begin
					state<=14;
					out<=50;
				end
				if(in == 517) begin
					state<=14;
					out<=51;
				end
				if(in == 518) begin
					state<=14;
					out<=52;
				end
				if(in == 519) begin
					state<=14;
					out<=53;
				end
				if(in == 520) begin
					state<=14;
					out<=54;
				end
				if(in == 521) begin
					state<=14;
					out<=55;
				end
				if(in == 522) begin
					state<=14;
					out<=56;
				end
				if(in == 523) begin
					state<=14;
					out<=57;
				end
				if(in == 524) begin
					state<=14;
					out<=58;
				end
				if(in == 525) begin
					state<=14;
					out<=59;
				end
				if(in == 526) begin
					state<=14;
					out<=60;
				end
				if(in == 527) begin
					state<=14;
					out<=61;
				end
				if(in == 528) begin
					state<=14;
					out<=62;
				end
				if(in == 529) begin
					state<=14;
					out<=63;
				end
				if(in == 530) begin
					state<=14;
					out<=64;
				end
				if(in == 531) begin
					state<=14;
					out<=65;
				end
				if(in == 532) begin
					state<=14;
					out<=66;
				end
				if(in == 533) begin
					state<=14;
					out<=67;
				end
				if(in == 534) begin
					state<=14;
					out<=68;
				end
				if(in == 535) begin
					state<=14;
					out<=69;
				end
				if(in == 536) begin
					state<=14;
					out<=70;
				end
				if(in == 537) begin
					state<=14;
					out<=71;
				end
				if(in == 538) begin
					state<=14;
					out<=72;
				end
				if(in == 539) begin
					state<=14;
					out<=73;
				end
				if(in == 540) begin
					state<=14;
					out<=74;
				end
				if(in == 541) begin
					state<=14;
					out<=75;
				end
				if(in == 542) begin
					state<=14;
					out<=76;
				end
				if(in == 543) begin
					state<=14;
					out<=77;
				end
				if(in == 544) begin
					state<=14;
					out<=78;
				end
				if(in == 545) begin
					state<=14;
					out<=79;
				end
				if(in == 546) begin
					state<=14;
					out<=80;
				end
				if(in == 547) begin
					state<=14;
					out<=81;
				end
				if(in == 548) begin
					state<=14;
					out<=82;
				end
				if(in == 549) begin
					state<=14;
					out<=83;
				end
				if(in == 550) begin
					state<=14;
					out<=84;
				end
				if(in == 551) begin
					state<=14;
					out<=85;
				end
				if(in == 552) begin
					state<=14;
					out<=86;
				end
				if(in == 553) begin
					state<=14;
					out<=87;
				end
				if(in == 554) begin
					state<=14;
					out<=88;
				end
				if(in == 555) begin
					state<=14;
					out<=89;
				end
				if(in == 556) begin
					state<=14;
					out<=90;
				end
				if(in == 557) begin
					state<=14;
					out<=91;
				end
				if(in == 558) begin
					state<=14;
					out<=92;
				end
				if(in == 559) begin
					state<=14;
					out<=93;
				end
				if(in == 560) begin
					state<=14;
					out<=94;
				end
				if(in == 561) begin
					state<=14;
					out<=95;
				end
				if(in == 562) begin
					state<=14;
					out<=96;
				end
				if(in == 563) begin
					state<=14;
					out<=97;
				end
				if(in == 564) begin
					state<=14;
					out<=98;
				end
				if(in == 565) begin
					state<=14;
					out<=99;
				end
				if(in == 566) begin
					state<=14;
					out<=100;
				end
				if(in == 567) begin
					state<=14;
					out<=101;
				end
				if(in == 568) begin
					state<=14;
					out<=102;
				end
				if(in == 569) begin
					state<=14;
					out<=103;
				end
				if(in == 570) begin
					state<=14;
					out<=104;
				end
				if(in == 571) begin
					state<=14;
					out<=105;
				end
				if(in == 572) begin
					state<=14;
					out<=106;
				end
				if(in == 573) begin
					state<=14;
					out<=107;
				end
				if(in == 574) begin
					state<=14;
					out<=108;
				end
				if(in == 575) begin
					state<=14;
					out<=109;
				end
				if(in == 576) begin
					state<=14;
					out<=110;
				end
				if(in == 577) begin
					state<=14;
					out<=111;
				end
				if(in == 578) begin
					state<=14;
					out<=112;
				end
				if(in == 579) begin
					state<=14;
					out<=113;
				end
				if(in == 580) begin
					state<=14;
					out<=114;
				end
				if(in == 581) begin
					state<=1;
					out<=115;
				end
				if(in == 582) begin
					state<=1;
					out<=116;
				end
				if(in == 583) begin
					state<=1;
					out<=117;
				end
				if(in == 584) begin
					state<=1;
					out<=118;
				end
				if(in == 585) begin
					state<=1;
					out<=119;
				end
				if(in == 586) begin
					state<=1;
					out<=120;
				end
				if(in == 587) begin
					state<=1;
					out<=121;
				end
				if(in == 588) begin
					state<=1;
					out<=122;
				end
				if(in == 589) begin
					state<=1;
					out<=123;
				end
				if(in == 590) begin
					state<=1;
					out<=124;
				end
				if(in == 591) begin
					state<=1;
					out<=125;
				end
				if(in == 592) begin
					state<=1;
					out<=126;
				end
				if(in == 593) begin
					state<=1;
					out<=127;
				end
				if(in == 594) begin
					state<=1;
					out<=128;
				end
				if(in == 595) begin
					state<=1;
					out<=129;
				end
				if(in == 596) begin
					state<=1;
					out<=130;
				end
				if(in == 597) begin
					state<=1;
					out<=131;
				end
				if(in == 598) begin
					state<=1;
					out<=132;
				end
				if(in == 599) begin
					state<=1;
					out<=133;
				end
				if(in == 600) begin
					state<=1;
					out<=134;
				end
				if(in == 601) begin
					state<=1;
					out<=135;
				end
				if(in == 602) begin
					state<=1;
					out<=136;
				end
				if(in == 603) begin
					state<=1;
					out<=137;
				end
				if(in == 604) begin
					state<=1;
					out<=138;
				end
				if(in == 605) begin
					state<=1;
					out<=139;
				end
				if(in == 606) begin
					state<=1;
					out<=140;
				end
				if(in == 607) begin
					state<=1;
					out<=141;
				end
				if(in == 608) begin
					state<=1;
					out<=142;
				end
				if(in == 609) begin
					state<=1;
					out<=143;
				end
				if(in == 610) begin
					state<=1;
					out<=144;
				end
				if(in == 611) begin
					state<=1;
					out<=145;
				end
				if(in == 612) begin
					state<=1;
					out<=146;
				end
				if(in == 613) begin
					state<=1;
					out<=147;
				end
				if(in == 614) begin
					state<=1;
					out<=148;
				end
				if(in == 615) begin
					state<=1;
					out<=149;
				end
				if(in == 616) begin
					state<=1;
					out<=150;
				end
				if(in == 617) begin
					state<=1;
					out<=151;
				end
				if(in == 618) begin
					state<=1;
					out<=152;
				end
				if(in == 619) begin
					state<=1;
					out<=153;
				end
				if(in == 620) begin
					state<=1;
					out<=154;
				end
				if(in == 621) begin
					state<=1;
					out<=155;
				end
				if(in == 622) begin
					state<=1;
					out<=156;
				end
				if(in == 623) begin
					state<=1;
					out<=157;
				end
				if(in == 624) begin
					state<=1;
					out<=158;
				end
				if(in == 625) begin
					state<=1;
					out<=159;
				end
				if(in == 626) begin
					state<=1;
					out<=160;
				end
				if(in == 627) begin
					state<=1;
					out<=161;
				end
				if(in == 628) begin
					state<=1;
					out<=162;
				end
				if(in == 629) begin
					state<=1;
					out<=163;
				end
				if(in == 630) begin
					state<=1;
					out<=164;
				end
				if(in == 631) begin
					state<=1;
					out<=165;
				end
				if(in == 632) begin
					state<=1;
					out<=166;
				end
				if(in == 633) begin
					state<=1;
					out<=167;
				end
				if(in == 634) begin
					state<=1;
					out<=168;
				end
				if(in == 635) begin
					state<=1;
					out<=169;
				end
				if(in == 636) begin
					state<=1;
					out<=170;
				end
				if(in == 637) begin
					state<=1;
					out<=171;
				end
				if(in == 638) begin
					state<=1;
					out<=172;
				end
				if(in == 639) begin
					state<=1;
					out<=173;
				end
				if(in == 640) begin
					state<=1;
					out<=174;
				end
				if(in == 641) begin
					state<=1;
					out<=175;
				end
				if(in == 642) begin
					state<=1;
					out<=176;
				end
				if(in == 643) begin
					state<=1;
					out<=177;
				end
				if(in == 644) begin
					state<=1;
					out<=178;
				end
				if(in == 645) begin
					state<=1;
					out<=179;
				end
				if(in == 646) begin
					state<=1;
					out<=180;
				end
				if(in == 647) begin
					state<=1;
					out<=181;
				end
				if(in == 648) begin
					state<=1;
					out<=182;
				end
				if(in == 649) begin
					state<=1;
					out<=183;
				end
				if(in == 650) begin
					state<=1;
					out<=184;
				end
				if(in == 651) begin
					state<=1;
					out<=185;
				end
				if(in == 652) begin
					state<=1;
					out<=186;
				end
				if(in == 653) begin
					state<=1;
					out<=187;
				end
				if(in == 654) begin
					state<=1;
					out<=188;
				end
				if(in == 655) begin
					state<=1;
					out<=189;
				end
				if(in == 656) begin
					state<=1;
					out<=190;
				end
				if(in == 657) begin
					state<=1;
					out<=191;
				end
				if(in == 658) begin
					state<=1;
					out<=192;
				end
				if(in == 659) begin
					state<=1;
					out<=193;
				end
				if(in == 660) begin
					state<=1;
					out<=194;
				end
				if(in == 661) begin
					state<=1;
					out<=195;
				end
				if(in == 662) begin
					state<=1;
					out<=196;
				end
				if(in == 663) begin
					state<=1;
					out<=197;
				end
				if(in == 664) begin
					state<=1;
					out<=198;
				end
				if(in == 665) begin
					state<=1;
					out<=199;
				end
				if(in == 666) begin
					state<=1;
					out<=200;
				end
				if(in == 667) begin
					state<=1;
					out<=201;
				end
				if(in == 668) begin
					state<=1;
					out<=202;
				end
				if(in == 669) begin
					state<=1;
					out<=203;
				end
				if(in == 670) begin
					state<=1;
					out<=204;
				end
				if(in == 671) begin
					state<=1;
					out<=205;
				end
				if(in == 672) begin
					state<=1;
					out<=206;
				end
				if(in == 673) begin
					state<=1;
					out<=207;
				end
				if(in == 674) begin
					state<=1;
					out<=208;
				end
				if(in == 675) begin
					state<=1;
					out<=209;
				end
				if(in == 676) begin
					state<=1;
					out<=210;
				end
				if(in == 677) begin
					state<=1;
					out<=211;
				end
				if(in == 678) begin
					state<=1;
					out<=212;
				end
				if(in == 679) begin
					state<=1;
					out<=213;
				end
				if(in == 680) begin
					state<=1;
					out<=214;
				end
				if(in == 681) begin
					state<=1;
					out<=215;
				end
				if(in == 682) begin
					state<=1;
					out<=216;
				end
				if(in == 683) begin
					state<=1;
					out<=217;
				end
				if(in == 684) begin
					state<=1;
					out<=218;
				end
				if(in == 685) begin
					state<=1;
					out<=219;
				end
				if(in == 686) begin
					state<=1;
					out<=220;
				end
				if(in == 687) begin
					state<=1;
					out<=221;
				end
				if(in == 688) begin
					state<=1;
					out<=222;
				end
				if(in == 689) begin
					state<=1;
					out<=223;
				end
				if(in == 690) begin
					state<=1;
					out<=224;
				end
				if(in == 691) begin
					state<=1;
					out<=225;
				end
				if(in == 692) begin
					state<=1;
					out<=226;
				end
				if(in == 693) begin
					state<=1;
					out<=227;
				end
				if(in == 694) begin
					state<=1;
					out<=228;
				end
				if(in == 695) begin
					state<=1;
					out<=229;
				end
				if(in == 696) begin
					state<=1;
					out<=230;
				end
				if(in == 697) begin
					state<=15;
					out<=231;
				end
				if(in == 698) begin
					state<=15;
					out<=232;
				end
				if(in == 699) begin
					state<=15;
					out<=233;
				end
				if(in == 700) begin
					state<=15;
					out<=234;
				end
				if(in == 701) begin
					state<=15;
					out<=235;
				end
				if(in == 702) begin
					state<=15;
					out<=236;
				end
				if(in == 703) begin
					state<=15;
					out<=237;
				end
				if(in == 704) begin
					state<=15;
					out<=238;
				end
				if(in == 705) begin
					state<=15;
					out<=239;
				end
				if(in == 706) begin
					state<=15;
					out<=240;
				end
				if(in == 707) begin
					state<=15;
					out<=241;
				end
				if(in == 708) begin
					state<=15;
					out<=242;
				end
				if(in == 709) begin
					state<=15;
					out<=243;
				end
				if(in == 710) begin
					state<=15;
					out<=244;
				end
				if(in == 711) begin
					state<=15;
					out<=245;
				end
				if(in == 712) begin
					state<=15;
					out<=246;
				end
				if(in == 713) begin
					state<=15;
					out<=247;
				end
				if(in == 714) begin
					state<=15;
					out<=248;
				end
				if(in == 715) begin
					state<=15;
					out<=249;
				end
				if(in == 716) begin
					state<=15;
					out<=250;
				end
				if(in == 717) begin
					state<=15;
					out<=251;
				end
				if(in == 718) begin
					state<=15;
					out<=252;
				end
				if(in == 719) begin
					state<=15;
					out<=253;
				end
				if(in == 720) begin
					state<=15;
					out<=254;
				end
				if(in == 721) begin
					state<=15;
					out<=255;
				end
				if(in == 722) begin
					state<=15;
					out<=0;
				end
				if(in == 723) begin
					state<=15;
					out<=1;
				end
				if(in == 724) begin
					state<=15;
					out<=2;
				end
				if(in == 725) begin
					state<=15;
					out<=3;
				end
				if(in == 726) begin
					state<=15;
					out<=4;
				end
				if(in == 727) begin
					state<=15;
					out<=5;
				end
				if(in == 728) begin
					state<=15;
					out<=6;
				end
				if(in == 729) begin
					state<=15;
					out<=7;
				end
				if(in == 730) begin
					state<=15;
					out<=8;
				end
				if(in == 731) begin
					state<=15;
					out<=9;
				end
				if(in == 732) begin
					state<=15;
					out<=10;
				end
				if(in == 733) begin
					state<=15;
					out<=11;
				end
				if(in == 734) begin
					state<=15;
					out<=12;
				end
				if(in == 735) begin
					state<=15;
					out<=13;
				end
				if(in == 736) begin
					state<=15;
					out<=14;
				end
				if(in == 737) begin
					state<=15;
					out<=15;
				end
				if(in == 738) begin
					state<=15;
					out<=16;
				end
				if(in == 739) begin
					state<=15;
					out<=17;
				end
				if(in == 740) begin
					state<=15;
					out<=18;
				end
				if(in == 741) begin
					state<=15;
					out<=19;
				end
				if(in == 742) begin
					state<=15;
					out<=20;
				end
				if(in == 743) begin
					state<=15;
					out<=21;
				end
				if(in == 744) begin
					state<=15;
					out<=22;
				end
				if(in == 745) begin
					state<=15;
					out<=23;
				end
				if(in == 746) begin
					state<=15;
					out<=24;
				end
				if(in == 747) begin
					state<=15;
					out<=25;
				end
				if(in == 748) begin
					state<=15;
					out<=26;
				end
				if(in == 749) begin
					state<=15;
					out<=27;
				end
				if(in == 750) begin
					state<=15;
					out<=28;
				end
				if(in == 751) begin
					state<=15;
					out<=29;
				end
				if(in == 752) begin
					state<=15;
					out<=30;
				end
				if(in == 753) begin
					state<=15;
					out<=31;
				end
				if(in == 754) begin
					state<=15;
					out<=32;
				end
				if(in == 755) begin
					state<=15;
					out<=33;
				end
				if(in == 756) begin
					state<=15;
					out<=34;
				end
				if(in == 757) begin
					state<=15;
					out<=35;
				end
				if(in == 758) begin
					state<=15;
					out<=36;
				end
				if(in == 759) begin
					state<=15;
					out<=37;
				end
				if(in == 760) begin
					state<=15;
					out<=38;
				end
				if(in == 761) begin
					state<=15;
					out<=39;
				end
				if(in == 762) begin
					state<=15;
					out<=40;
				end
				if(in == 763) begin
					state<=15;
					out<=41;
				end
				if(in == 764) begin
					state<=15;
					out<=42;
				end
				if(in == 765) begin
					state<=15;
					out<=43;
				end
				if(in == 766) begin
					state<=15;
					out<=44;
				end
				if(in == 767) begin
					state<=15;
					out<=45;
				end
				if(in == 768) begin
					state<=15;
					out<=46;
				end
				if(in == 769) begin
					state<=15;
					out<=47;
				end
				if(in == 770) begin
					state<=15;
					out<=48;
				end
				if(in == 771) begin
					state<=15;
					out<=49;
				end
				if(in == 772) begin
					state<=15;
					out<=50;
				end
				if(in == 773) begin
					state<=15;
					out<=51;
				end
				if(in == 774) begin
					state<=15;
					out<=52;
				end
				if(in == 775) begin
					state<=15;
					out<=53;
				end
				if(in == 776) begin
					state<=15;
					out<=54;
				end
				if(in == 777) begin
					state<=15;
					out<=55;
				end
				if(in == 778) begin
					state<=15;
					out<=56;
				end
				if(in == 779) begin
					state<=15;
					out<=57;
				end
				if(in == 780) begin
					state<=15;
					out<=58;
				end
				if(in == 781) begin
					state<=15;
					out<=59;
				end
				if(in == 782) begin
					state<=15;
					out<=60;
				end
				if(in == 783) begin
					state<=15;
					out<=61;
				end
				if(in == 784) begin
					state<=15;
					out<=62;
				end
				if(in == 785) begin
					state<=15;
					out<=63;
				end
				if(in == 786) begin
					state<=15;
					out<=64;
				end
				if(in == 787) begin
					state<=15;
					out<=65;
				end
				if(in == 788) begin
					state<=15;
					out<=66;
				end
				if(in == 789) begin
					state<=15;
					out<=67;
				end
				if(in == 790) begin
					state<=15;
					out<=68;
				end
				if(in == 791) begin
					state<=15;
					out<=69;
				end
				if(in == 792) begin
					state<=15;
					out<=70;
				end
				if(in == 793) begin
					state<=15;
					out<=71;
				end
				if(in == 794) begin
					state<=15;
					out<=72;
				end
				if(in == 795) begin
					state<=15;
					out<=73;
				end
				if(in == 796) begin
					state<=15;
					out<=74;
				end
				if(in == 797) begin
					state<=15;
					out<=75;
				end
				if(in == 798) begin
					state<=15;
					out<=76;
				end
				if(in == 799) begin
					state<=15;
					out<=77;
				end
				if(in == 800) begin
					state<=15;
					out<=78;
				end
				if(in == 801) begin
					state<=15;
					out<=79;
				end
				if(in == 802) begin
					state<=15;
					out<=80;
				end
				if(in == 803) begin
					state<=15;
					out<=81;
				end
				if(in == 804) begin
					state<=15;
					out<=82;
				end
				if(in == 805) begin
					state<=15;
					out<=83;
				end
				if(in == 806) begin
					state<=15;
					out<=84;
				end
				if(in == 807) begin
					state<=15;
					out<=85;
				end
				if(in == 808) begin
					state<=15;
					out<=86;
				end
				if(in == 809) begin
					state<=15;
					out<=87;
				end
				if(in == 810) begin
					state<=15;
					out<=88;
				end
				if(in == 811) begin
					state<=15;
					out<=89;
				end
				if(in == 812) begin
					state<=15;
					out<=90;
				end
				if(in == 813) begin
					state<=16;
					out<=91;
				end
				if(in == 814) begin
					state<=16;
					out<=92;
				end
				if(in == 815) begin
					state<=16;
					out<=93;
				end
				if(in == 816) begin
					state<=16;
					out<=94;
				end
				if(in == 817) begin
					state<=16;
					out<=95;
				end
				if(in == 818) begin
					state<=16;
					out<=96;
				end
				if(in == 819) begin
					state<=16;
					out<=97;
				end
				if(in == 820) begin
					state<=16;
					out<=98;
				end
				if(in == 821) begin
					state<=16;
					out<=99;
				end
				if(in == 822) begin
					state<=16;
					out<=100;
				end
				if(in == 823) begin
					state<=16;
					out<=101;
				end
				if(in == 824) begin
					state<=16;
					out<=102;
				end
				if(in == 825) begin
					state<=16;
					out<=103;
				end
				if(in == 826) begin
					state<=16;
					out<=104;
				end
				if(in == 827) begin
					state<=16;
					out<=105;
				end
				if(in == 828) begin
					state<=16;
					out<=106;
				end
				if(in == 829) begin
					state<=16;
					out<=107;
				end
				if(in == 830) begin
					state<=16;
					out<=108;
				end
				if(in == 831) begin
					state<=16;
					out<=109;
				end
				if(in == 832) begin
					state<=16;
					out<=110;
				end
				if(in == 833) begin
					state<=16;
					out<=111;
				end
				if(in == 834) begin
					state<=16;
					out<=112;
				end
				if(in == 835) begin
					state<=16;
					out<=113;
				end
				if(in == 836) begin
					state<=16;
					out<=114;
				end
				if(in == 837) begin
					state<=16;
					out<=115;
				end
				if(in == 838) begin
					state<=16;
					out<=116;
				end
				if(in == 839) begin
					state<=16;
					out<=117;
				end
				if(in == 840) begin
					state<=16;
					out<=118;
				end
				if(in == 841) begin
					state<=16;
					out<=119;
				end
				if(in == 842) begin
					state<=16;
					out<=120;
				end
				if(in == 843) begin
					state<=16;
					out<=121;
				end
				if(in == 844) begin
					state<=16;
					out<=122;
				end
				if(in == 845) begin
					state<=16;
					out<=123;
				end
				if(in == 846) begin
					state<=16;
					out<=124;
				end
				if(in == 847) begin
					state<=16;
					out<=125;
				end
				if(in == 848) begin
					state<=16;
					out<=126;
				end
				if(in == 849) begin
					state<=16;
					out<=127;
				end
				if(in == 850) begin
					state<=16;
					out<=128;
				end
				if(in == 851) begin
					state<=16;
					out<=129;
				end
				if(in == 852) begin
					state<=16;
					out<=130;
				end
				if(in == 853) begin
					state<=16;
					out<=131;
				end
				if(in == 854) begin
					state<=16;
					out<=132;
				end
				if(in == 855) begin
					state<=16;
					out<=133;
				end
				if(in == 856) begin
					state<=16;
					out<=134;
				end
				if(in == 857) begin
					state<=16;
					out<=135;
				end
				if(in == 858) begin
					state<=16;
					out<=136;
				end
				if(in == 859) begin
					state<=16;
					out<=137;
				end
				if(in == 860) begin
					state<=16;
					out<=138;
				end
				if(in == 861) begin
					state<=16;
					out<=139;
				end
				if(in == 862) begin
					state<=16;
					out<=140;
				end
				if(in == 863) begin
					state<=16;
					out<=141;
				end
				if(in == 864) begin
					state<=16;
					out<=142;
				end
				if(in == 865) begin
					state<=16;
					out<=143;
				end
				if(in == 866) begin
					state<=16;
					out<=144;
				end
				if(in == 867) begin
					state<=16;
					out<=145;
				end
				if(in == 868) begin
					state<=16;
					out<=146;
				end
				if(in == 869) begin
					state<=16;
					out<=147;
				end
				if(in == 870) begin
					state<=16;
					out<=148;
				end
				if(in == 871) begin
					state<=16;
					out<=149;
				end
				if(in == 872) begin
					state<=16;
					out<=150;
				end
				if(in == 873) begin
					state<=16;
					out<=151;
				end
				if(in == 874) begin
					state<=16;
					out<=152;
				end
				if(in == 875) begin
					state<=16;
					out<=153;
				end
				if(in == 876) begin
					state<=16;
					out<=154;
				end
				if(in == 877) begin
					state<=16;
					out<=155;
				end
				if(in == 878) begin
					state<=16;
					out<=156;
				end
				if(in == 879) begin
					state<=16;
					out<=157;
				end
				if(in == 880) begin
					state<=16;
					out<=158;
				end
				if(in == 881) begin
					state<=16;
					out<=159;
				end
				if(in == 882) begin
					state<=16;
					out<=160;
				end
				if(in == 883) begin
					state<=16;
					out<=161;
				end
				if(in == 884) begin
					state<=16;
					out<=162;
				end
				if(in == 885) begin
					state<=16;
					out<=163;
				end
				if(in == 886) begin
					state<=16;
					out<=164;
				end
				if(in == 887) begin
					state<=16;
					out<=165;
				end
				if(in == 888) begin
					state<=16;
					out<=166;
				end
				if(in == 889) begin
					state<=16;
					out<=167;
				end
				if(in == 890) begin
					state<=16;
					out<=168;
				end
				if(in == 891) begin
					state<=16;
					out<=169;
				end
				if(in == 892) begin
					state<=16;
					out<=170;
				end
				if(in == 893) begin
					state<=16;
					out<=171;
				end
				if(in == 894) begin
					state<=16;
					out<=172;
				end
				if(in == 895) begin
					state<=16;
					out<=173;
				end
				if(in == 896) begin
					state<=16;
					out<=174;
				end
				if(in == 897) begin
					state<=16;
					out<=175;
				end
				if(in == 898) begin
					state<=16;
					out<=176;
				end
				if(in == 899) begin
					state<=16;
					out<=177;
				end
				if(in == 900) begin
					state<=16;
					out<=178;
				end
				if(in == 901) begin
					state<=16;
					out<=179;
				end
				if(in == 902) begin
					state<=16;
					out<=180;
				end
				if(in == 903) begin
					state<=16;
					out<=181;
				end
				if(in == 904) begin
					state<=16;
					out<=182;
				end
				if(in == 905) begin
					state<=16;
					out<=183;
				end
				if(in == 906) begin
					state<=16;
					out<=184;
				end
				if(in == 907) begin
					state<=16;
					out<=185;
				end
				if(in == 908) begin
					state<=16;
					out<=186;
				end
				if(in == 909) begin
					state<=16;
					out<=187;
				end
				if(in == 910) begin
					state<=16;
					out<=188;
				end
				if(in == 911) begin
					state<=16;
					out<=189;
				end
				if(in == 912) begin
					state<=16;
					out<=190;
				end
				if(in == 913) begin
					state<=16;
					out<=191;
				end
				if(in == 914) begin
					state<=16;
					out<=192;
				end
				if(in == 915) begin
					state<=16;
					out<=193;
				end
				if(in == 916) begin
					state<=16;
					out<=194;
				end
				if(in == 917) begin
					state<=16;
					out<=195;
				end
				if(in == 918) begin
					state<=16;
					out<=196;
				end
				if(in == 919) begin
					state<=16;
					out<=197;
				end
				if(in == 920) begin
					state<=16;
					out<=198;
				end
				if(in == 921) begin
					state<=16;
					out<=199;
				end
				if(in == 922) begin
					state<=16;
					out<=200;
				end
				if(in == 923) begin
					state<=16;
					out<=201;
				end
				if(in == 924) begin
					state<=16;
					out<=202;
				end
				if(in == 925) begin
					state<=16;
					out<=203;
				end
				if(in == 926) begin
					state<=16;
					out<=204;
				end
				if(in == 927) begin
					state<=16;
					out<=205;
				end
				if(in == 928) begin
					state<=16;
					out<=206;
				end
			end
			15: begin
				if(in == 0) begin
					state<=2;
					out<=207;
				end
				if(in == 1) begin
					state<=1;
					out<=208;
				end
				if(in == 2) begin
					state<=2;
					out<=209;
				end
				if(in == 3) begin
					state<=2;
					out<=210;
				end
				if(in == 4) begin
					state<=2;
					out<=211;
				end
				if(in == 5) begin
					state<=2;
					out<=212;
				end
				if(in == 6) begin
					state<=2;
					out<=213;
				end
				if(in == 7) begin
					state<=2;
					out<=214;
				end
				if(in == 8) begin
					state<=2;
					out<=215;
				end
				if(in == 9) begin
					state<=2;
					out<=216;
				end
				if(in == 10) begin
					state<=2;
					out<=217;
				end
				if(in == 11) begin
					state<=2;
					out<=218;
				end
				if(in == 12) begin
					state<=2;
					out<=219;
				end
				if(in == 13) begin
					state<=2;
					out<=220;
				end
				if(in == 14) begin
					state<=2;
					out<=221;
				end
				if(in == 15) begin
					state<=2;
					out<=222;
				end
				if(in == 16) begin
					state<=2;
					out<=223;
				end
				if(in == 17) begin
					state<=2;
					out<=224;
				end
				if(in == 18) begin
					state<=2;
					out<=225;
				end
				if(in == 19) begin
					state<=2;
					out<=226;
				end
				if(in == 20) begin
					state<=2;
					out<=227;
				end
				if(in == 21) begin
					state<=2;
					out<=228;
				end
				if(in == 22) begin
					state<=2;
					out<=229;
				end
				if(in == 23) begin
					state<=2;
					out<=230;
				end
				if(in == 24) begin
					state<=2;
					out<=231;
				end
				if(in == 25) begin
					state<=2;
					out<=232;
				end
				if(in == 26) begin
					state<=2;
					out<=233;
				end
				if(in == 27) begin
					state<=2;
					out<=234;
				end
				if(in == 28) begin
					state<=2;
					out<=235;
				end
				if(in == 29) begin
					state<=2;
					out<=236;
				end
				if(in == 30) begin
					state<=2;
					out<=237;
				end
				if(in == 31) begin
					state<=2;
					out<=238;
				end
				if(in == 32) begin
					state<=2;
					out<=239;
				end
				if(in == 33) begin
					state<=2;
					out<=240;
				end
				if(in == 34) begin
					state<=2;
					out<=241;
				end
				if(in == 35) begin
					state<=2;
					out<=242;
				end
				if(in == 36) begin
					state<=2;
					out<=243;
				end
				if(in == 37) begin
					state<=2;
					out<=244;
				end
				if(in == 38) begin
					state<=2;
					out<=245;
				end
				if(in == 39) begin
					state<=2;
					out<=246;
				end
				if(in == 40) begin
					state<=2;
					out<=247;
				end
				if(in == 41) begin
					state<=2;
					out<=248;
				end
				if(in == 42) begin
					state<=2;
					out<=249;
				end
				if(in == 43) begin
					state<=2;
					out<=250;
				end
				if(in == 44) begin
					state<=2;
					out<=251;
				end
				if(in == 45) begin
					state<=2;
					out<=252;
				end
				if(in == 46) begin
					state<=2;
					out<=253;
				end
				if(in == 47) begin
					state<=2;
					out<=254;
				end
				if(in == 48) begin
					state<=2;
					out<=255;
				end
				if(in == 49) begin
					state<=2;
					out<=0;
				end
				if(in == 50) begin
					state<=2;
					out<=1;
				end
				if(in == 51) begin
					state<=2;
					out<=2;
				end
				if(in == 52) begin
					state<=2;
					out<=3;
				end
				if(in == 53) begin
					state<=2;
					out<=4;
				end
				if(in == 54) begin
					state<=2;
					out<=5;
				end
				if(in == 55) begin
					state<=2;
					out<=6;
				end
				if(in == 56) begin
					state<=2;
					out<=7;
				end
				if(in == 57) begin
					state<=2;
					out<=8;
				end
				if(in == 58) begin
					state<=2;
					out<=9;
				end
				if(in == 59) begin
					state<=2;
					out<=10;
				end
				if(in == 60) begin
					state<=2;
					out<=11;
				end
				if(in == 61) begin
					state<=2;
					out<=12;
				end
				if(in == 62) begin
					state<=2;
					out<=13;
				end
				if(in == 63) begin
					state<=2;
					out<=14;
				end
				if(in == 64) begin
					state<=2;
					out<=15;
				end
				if(in == 65) begin
					state<=2;
					out<=16;
				end
				if(in == 66) begin
					state<=2;
					out<=17;
				end
				if(in == 67) begin
					state<=2;
					out<=18;
				end
				if(in == 68) begin
					state<=2;
					out<=19;
				end
				if(in == 69) begin
					state<=2;
					out<=20;
				end
				if(in == 70) begin
					state<=2;
					out<=21;
				end
				if(in == 71) begin
					state<=2;
					out<=22;
				end
				if(in == 72) begin
					state<=2;
					out<=23;
				end
				if(in == 73) begin
					state<=2;
					out<=24;
				end
				if(in == 74) begin
					state<=2;
					out<=25;
				end
				if(in == 75) begin
					state<=2;
					out<=26;
				end
				if(in == 76) begin
					state<=2;
					out<=27;
				end
				if(in == 77) begin
					state<=2;
					out<=28;
				end
				if(in == 78) begin
					state<=2;
					out<=29;
				end
				if(in == 79) begin
					state<=2;
					out<=30;
				end
				if(in == 80) begin
					state<=2;
					out<=31;
				end
				if(in == 81) begin
					state<=2;
					out<=32;
				end
				if(in == 82) begin
					state<=2;
					out<=33;
				end
				if(in == 83) begin
					state<=2;
					out<=34;
				end
				if(in == 84) begin
					state<=2;
					out<=35;
				end
				if(in == 85) begin
					state<=2;
					out<=36;
				end
				if(in == 86) begin
					state<=2;
					out<=37;
				end
				if(in == 87) begin
					state<=2;
					out<=38;
				end
				if(in == 88) begin
					state<=2;
					out<=39;
				end
				if(in == 89) begin
					state<=2;
					out<=40;
				end
				if(in == 90) begin
					state<=2;
					out<=41;
				end
				if(in == 91) begin
					state<=2;
					out<=42;
				end
				if(in == 92) begin
					state<=2;
					out<=43;
				end
				if(in == 93) begin
					state<=2;
					out<=44;
				end
				if(in == 94) begin
					state<=2;
					out<=45;
				end
				if(in == 95) begin
					state<=2;
					out<=46;
				end
				if(in == 96) begin
					state<=2;
					out<=47;
				end
				if(in == 97) begin
					state<=2;
					out<=48;
				end
				if(in == 98) begin
					state<=2;
					out<=49;
				end
				if(in == 99) begin
					state<=2;
					out<=50;
				end
				if(in == 100) begin
					state<=2;
					out<=51;
				end
				if(in == 101) begin
					state<=2;
					out<=52;
				end
				if(in == 102) begin
					state<=2;
					out<=53;
				end
				if(in == 103) begin
					state<=2;
					out<=54;
				end
				if(in == 104) begin
					state<=2;
					out<=55;
				end
				if(in == 105) begin
					state<=2;
					out<=56;
				end
				if(in == 106) begin
					state<=2;
					out<=57;
				end
				if(in == 107) begin
					state<=2;
					out<=58;
				end
				if(in == 108) begin
					state<=2;
					out<=59;
				end
				if(in == 109) begin
					state<=2;
					out<=60;
				end
				if(in == 110) begin
					state<=2;
					out<=61;
				end
				if(in == 111) begin
					state<=2;
					out<=62;
				end
				if(in == 112) begin
					state<=2;
					out<=63;
				end
				if(in == 113) begin
					state<=2;
					out<=64;
				end
				if(in == 114) begin
					state<=2;
					out<=65;
				end
				if(in == 115) begin
					state<=2;
					out<=66;
				end
				if(in == 116) begin
					state<=2;
					out<=67;
				end
				if(in == 117) begin
					state<=2;
					out<=68;
				end
				if(in == 118) begin
					state<=2;
					out<=69;
				end
				if(in == 119) begin
					state<=2;
					out<=70;
				end
				if(in == 120) begin
					state<=2;
					out<=71;
				end
				if(in == 121) begin
					state<=2;
					out<=72;
				end
				if(in == 122) begin
					state<=2;
					out<=73;
				end
				if(in == 123) begin
					state<=2;
					out<=74;
				end
				if(in == 124) begin
					state<=2;
					out<=75;
				end
				if(in == 125) begin
					state<=2;
					out<=76;
				end
				if(in == 126) begin
					state<=2;
					out<=77;
				end
				if(in == 127) begin
					state<=2;
					out<=78;
				end
				if(in == 128) begin
					state<=2;
					out<=79;
				end
				if(in == 129) begin
					state<=2;
					out<=80;
				end
				if(in == 130) begin
					state<=2;
					out<=81;
				end
				if(in == 131) begin
					state<=2;
					out<=82;
				end
				if(in == 132) begin
					state<=2;
					out<=83;
				end
				if(in == 133) begin
					state<=2;
					out<=84;
				end
				if(in == 134) begin
					state<=2;
					out<=85;
				end
				if(in == 135) begin
					state<=2;
					out<=86;
				end
				if(in == 136) begin
					state<=2;
					out<=87;
				end
				if(in == 137) begin
					state<=2;
					out<=88;
				end
				if(in == 138) begin
					state<=2;
					out<=89;
				end
				if(in == 139) begin
					state<=2;
					out<=90;
				end
				if(in == 140) begin
					state<=2;
					out<=91;
				end
				if(in == 141) begin
					state<=2;
					out<=92;
				end
				if(in == 142) begin
					state<=2;
					out<=93;
				end
				if(in == 143) begin
					state<=2;
					out<=94;
				end
				if(in == 144) begin
					state<=2;
					out<=95;
				end
				if(in == 145) begin
					state<=2;
					out<=96;
				end
				if(in == 146) begin
					state<=2;
					out<=97;
				end
				if(in == 147) begin
					state<=2;
					out<=98;
				end
				if(in == 148) begin
					state<=2;
					out<=99;
				end
				if(in == 149) begin
					state<=2;
					out<=100;
				end
				if(in == 150) begin
					state<=2;
					out<=101;
				end
				if(in == 151) begin
					state<=2;
					out<=102;
				end
				if(in == 152) begin
					state<=2;
					out<=103;
				end
				if(in == 153) begin
					state<=2;
					out<=104;
				end
				if(in == 154) begin
					state<=2;
					out<=105;
				end
				if(in == 155) begin
					state<=2;
					out<=106;
				end
				if(in == 156) begin
					state<=2;
					out<=107;
				end
				if(in == 157) begin
					state<=2;
					out<=108;
				end
				if(in == 158) begin
					state<=2;
					out<=109;
				end
				if(in == 159) begin
					state<=2;
					out<=110;
				end
				if(in == 160) begin
					state<=2;
					out<=111;
				end
				if(in == 161) begin
					state<=2;
					out<=112;
				end
				if(in == 162) begin
					state<=2;
					out<=113;
				end
				if(in == 163) begin
					state<=2;
					out<=114;
				end
				if(in == 164) begin
					state<=2;
					out<=115;
				end
				if(in == 165) begin
					state<=2;
					out<=116;
				end
				if(in == 166) begin
					state<=2;
					out<=117;
				end
				if(in == 167) begin
					state<=2;
					out<=118;
				end
				if(in == 168) begin
					state<=2;
					out<=119;
				end
				if(in == 169) begin
					state<=2;
					out<=120;
				end
				if(in == 170) begin
					state<=2;
					out<=121;
				end
				if(in == 171) begin
					state<=2;
					out<=122;
				end
				if(in == 172) begin
					state<=2;
					out<=123;
				end
				if(in == 173) begin
					state<=2;
					out<=124;
				end
				if(in == 174) begin
					state<=2;
					out<=125;
				end
				if(in == 175) begin
					state<=2;
					out<=126;
				end
				if(in == 176) begin
					state<=2;
					out<=127;
				end
				if(in == 177) begin
					state<=2;
					out<=128;
				end
				if(in == 178) begin
					state<=2;
					out<=129;
				end
				if(in == 179) begin
					state<=2;
					out<=130;
				end
				if(in == 180) begin
					state<=2;
					out<=131;
				end
				if(in == 181) begin
					state<=2;
					out<=132;
				end
				if(in == 182) begin
					state<=2;
					out<=133;
				end
				if(in == 183) begin
					state<=2;
					out<=134;
				end
				if(in == 184) begin
					state<=2;
					out<=135;
				end
				if(in == 185) begin
					state<=2;
					out<=136;
				end
				if(in == 186) begin
					state<=2;
					out<=137;
				end
				if(in == 187) begin
					state<=2;
					out<=138;
				end
				if(in == 188) begin
					state<=2;
					out<=139;
				end
				if(in == 189) begin
					state<=2;
					out<=140;
				end
				if(in == 190) begin
					state<=2;
					out<=141;
				end
				if(in == 191) begin
					state<=2;
					out<=142;
				end
				if(in == 192) begin
					state<=2;
					out<=143;
				end
				if(in == 193) begin
					state<=2;
					out<=144;
				end
				if(in == 194) begin
					state<=2;
					out<=145;
				end
				if(in == 195) begin
					state<=2;
					out<=146;
				end
				if(in == 196) begin
					state<=2;
					out<=147;
				end
				if(in == 197) begin
					state<=2;
					out<=148;
				end
				if(in == 198) begin
					state<=2;
					out<=149;
				end
				if(in == 199) begin
					state<=2;
					out<=150;
				end
				if(in == 200) begin
					state<=2;
					out<=151;
				end
				if(in == 201) begin
					state<=2;
					out<=152;
				end
				if(in == 202) begin
					state<=2;
					out<=153;
				end
				if(in == 203) begin
					state<=2;
					out<=154;
				end
				if(in == 204) begin
					state<=2;
					out<=155;
				end
				if(in == 205) begin
					state<=2;
					out<=156;
				end
				if(in == 206) begin
					state<=2;
					out<=157;
				end
				if(in == 207) begin
					state<=2;
					out<=158;
				end
				if(in == 208) begin
					state<=2;
					out<=159;
				end
				if(in == 209) begin
					state<=2;
					out<=160;
				end
				if(in == 210) begin
					state<=2;
					out<=161;
				end
				if(in == 211) begin
					state<=2;
					out<=162;
				end
				if(in == 212) begin
					state<=2;
					out<=163;
				end
				if(in == 213) begin
					state<=2;
					out<=164;
				end
				if(in == 214) begin
					state<=2;
					out<=165;
				end
				if(in == 215) begin
					state<=2;
					out<=166;
				end
				if(in == 216) begin
					state<=2;
					out<=167;
				end
				if(in == 217) begin
					state<=2;
					out<=168;
				end
				if(in == 218) begin
					state<=2;
					out<=169;
				end
				if(in == 219) begin
					state<=2;
					out<=170;
				end
				if(in == 220) begin
					state<=2;
					out<=171;
				end
				if(in == 221) begin
					state<=2;
					out<=172;
				end
				if(in == 222) begin
					state<=2;
					out<=173;
				end
				if(in == 223) begin
					state<=2;
					out<=174;
				end
				if(in == 224) begin
					state<=2;
					out<=175;
				end
				if(in == 225) begin
					state<=2;
					out<=176;
				end
				if(in == 226) begin
					state<=2;
					out<=177;
				end
				if(in == 227) begin
					state<=2;
					out<=178;
				end
				if(in == 228) begin
					state<=2;
					out<=179;
				end
				if(in == 229) begin
					state<=2;
					out<=180;
				end
				if(in == 230) begin
					state<=2;
					out<=181;
				end
				if(in == 231) begin
					state<=2;
					out<=182;
				end
				if(in == 232) begin
					state<=2;
					out<=183;
				end
				if(in == 233) begin
					state<=2;
					out<=184;
				end
				if(in == 234) begin
					state<=2;
					out<=185;
				end
				if(in == 235) begin
					state<=2;
					out<=186;
				end
				if(in == 236) begin
					state<=2;
					out<=187;
				end
				if(in == 237) begin
					state<=2;
					out<=188;
				end
				if(in == 238) begin
					state<=2;
					out<=189;
				end
				if(in == 239) begin
					state<=2;
					out<=190;
				end
				if(in == 240) begin
					state<=2;
					out<=191;
				end
				if(in == 241) begin
					state<=2;
					out<=192;
				end
				if(in == 242) begin
					state<=2;
					out<=193;
				end
				if(in == 243) begin
					state<=2;
					out<=194;
				end
				if(in == 244) begin
					state<=2;
					out<=195;
				end
				if(in == 245) begin
					state<=2;
					out<=196;
				end
				if(in == 246) begin
					state<=2;
					out<=197;
				end
				if(in == 247) begin
					state<=2;
					out<=198;
				end
				if(in == 248) begin
					state<=2;
					out<=199;
				end
				if(in == 249) begin
					state<=2;
					out<=200;
				end
				if(in == 250) begin
					state<=2;
					out<=201;
				end
				if(in == 251) begin
					state<=2;
					out<=202;
				end
				if(in == 252) begin
					state<=2;
					out<=203;
				end
				if(in == 253) begin
					state<=2;
					out<=204;
				end
				if(in == 254) begin
					state<=2;
					out<=205;
				end
				if(in == 255) begin
					state<=2;
					out<=206;
				end
				if(in == 256) begin
					state<=2;
					out<=207;
				end
				if(in == 257) begin
					state<=2;
					out<=208;
				end
				if(in == 258) begin
					state<=2;
					out<=209;
				end
				if(in == 259) begin
					state<=2;
					out<=210;
				end
				if(in == 260) begin
					state<=2;
					out<=211;
				end
				if(in == 261) begin
					state<=2;
					out<=212;
				end
				if(in == 262) begin
					state<=2;
					out<=213;
				end
				if(in == 263) begin
					state<=2;
					out<=214;
				end
				if(in == 264) begin
					state<=2;
					out<=215;
				end
				if(in == 265) begin
					state<=2;
					out<=216;
				end
				if(in == 266) begin
					state<=2;
					out<=217;
				end
				if(in == 267) begin
					state<=2;
					out<=218;
				end
				if(in == 268) begin
					state<=2;
					out<=219;
				end
				if(in == 269) begin
					state<=2;
					out<=220;
				end
				if(in == 270) begin
					state<=2;
					out<=221;
				end
				if(in == 271) begin
					state<=2;
					out<=222;
				end
				if(in == 272) begin
					state<=2;
					out<=223;
				end
				if(in == 273) begin
					state<=2;
					out<=224;
				end
				if(in == 274) begin
					state<=2;
					out<=225;
				end
				if(in == 275) begin
					state<=2;
					out<=226;
				end
				if(in == 276) begin
					state<=2;
					out<=227;
				end
				if(in == 277) begin
					state<=2;
					out<=228;
				end
				if(in == 278) begin
					state<=2;
					out<=229;
				end
				if(in == 279) begin
					state<=2;
					out<=230;
				end
				if(in == 280) begin
					state<=2;
					out<=231;
				end
				if(in == 281) begin
					state<=2;
					out<=232;
				end
				if(in == 282) begin
					state<=2;
					out<=233;
				end
				if(in == 283) begin
					state<=2;
					out<=234;
				end
				if(in == 284) begin
					state<=2;
					out<=235;
				end
				if(in == 285) begin
					state<=2;
					out<=236;
				end
				if(in == 286) begin
					state<=2;
					out<=237;
				end
				if(in == 287) begin
					state<=2;
					out<=238;
				end
				if(in == 288) begin
					state<=2;
					out<=239;
				end
				if(in == 289) begin
					state<=2;
					out<=240;
				end
				if(in == 290) begin
					state<=2;
					out<=241;
				end
				if(in == 291) begin
					state<=2;
					out<=242;
				end
				if(in == 292) begin
					state<=2;
					out<=243;
				end
				if(in == 293) begin
					state<=2;
					out<=244;
				end
				if(in == 294) begin
					state<=2;
					out<=245;
				end
				if(in == 295) begin
					state<=2;
					out<=246;
				end
				if(in == 296) begin
					state<=2;
					out<=247;
				end
				if(in == 297) begin
					state<=2;
					out<=248;
				end
				if(in == 298) begin
					state<=2;
					out<=249;
				end
				if(in == 299) begin
					state<=2;
					out<=250;
				end
				if(in == 300) begin
					state<=2;
					out<=251;
				end
				if(in == 301) begin
					state<=2;
					out<=252;
				end
				if(in == 302) begin
					state<=2;
					out<=253;
				end
				if(in == 303) begin
					state<=2;
					out<=254;
				end
				if(in == 304) begin
					state<=2;
					out<=255;
				end
				if(in == 305) begin
					state<=2;
					out<=0;
				end
				if(in == 306) begin
					state<=2;
					out<=1;
				end
				if(in == 307) begin
					state<=2;
					out<=2;
				end
				if(in == 308) begin
					state<=2;
					out<=3;
				end
				if(in == 309) begin
					state<=2;
					out<=4;
				end
				if(in == 310) begin
					state<=2;
					out<=5;
				end
				if(in == 311) begin
					state<=2;
					out<=6;
				end
				if(in == 312) begin
					state<=2;
					out<=7;
				end
				if(in == 313) begin
					state<=2;
					out<=8;
				end
				if(in == 314) begin
					state<=2;
					out<=9;
				end
				if(in == 315) begin
					state<=2;
					out<=10;
				end
				if(in == 316) begin
					state<=2;
					out<=11;
				end
				if(in == 317) begin
					state<=2;
					out<=12;
				end
				if(in == 318) begin
					state<=2;
					out<=13;
				end
				if(in == 319) begin
					state<=2;
					out<=14;
				end
				if(in == 320) begin
					state<=2;
					out<=15;
				end
				if(in == 321) begin
					state<=2;
					out<=16;
				end
				if(in == 322) begin
					state<=2;
					out<=17;
				end
				if(in == 323) begin
					state<=2;
					out<=18;
				end
				if(in == 324) begin
					state<=2;
					out<=19;
				end
				if(in == 325) begin
					state<=2;
					out<=20;
				end
				if(in == 326) begin
					state<=2;
					out<=21;
				end
				if(in == 327) begin
					state<=2;
					out<=22;
				end
				if(in == 328) begin
					state<=2;
					out<=23;
				end
				if(in == 329) begin
					state<=2;
					out<=24;
				end
				if(in == 330) begin
					state<=2;
					out<=25;
				end
				if(in == 331) begin
					state<=2;
					out<=26;
				end
				if(in == 332) begin
					state<=2;
					out<=27;
				end
				if(in == 333) begin
					state<=2;
					out<=28;
				end
				if(in == 334) begin
					state<=2;
					out<=29;
				end
				if(in == 335) begin
					state<=2;
					out<=30;
				end
				if(in == 336) begin
					state<=2;
					out<=31;
				end
				if(in == 337) begin
					state<=2;
					out<=32;
				end
				if(in == 338) begin
					state<=2;
					out<=33;
				end
				if(in == 339) begin
					state<=2;
					out<=34;
				end
				if(in == 340) begin
					state<=2;
					out<=35;
				end
				if(in == 341) begin
					state<=2;
					out<=36;
				end
				if(in == 342) begin
					state<=2;
					out<=37;
				end
				if(in == 343) begin
					state<=2;
					out<=38;
				end
				if(in == 344) begin
					state<=2;
					out<=39;
				end
				if(in == 345) begin
					state<=2;
					out<=40;
				end
				if(in == 346) begin
					state<=2;
					out<=41;
				end
				if(in == 347) begin
					state<=2;
					out<=42;
				end
				if(in == 348) begin
					state<=2;
					out<=43;
				end
				if(in == 349) begin
					state<=2;
					out<=44;
				end
				if(in == 350) begin
					state<=2;
					out<=45;
				end
				if(in == 351) begin
					state<=2;
					out<=46;
				end
				if(in == 352) begin
					state<=2;
					out<=47;
				end
				if(in == 353) begin
					state<=2;
					out<=48;
				end
				if(in == 354) begin
					state<=2;
					out<=49;
				end
				if(in == 355) begin
					state<=2;
					out<=50;
				end
				if(in == 356) begin
					state<=2;
					out<=51;
				end
				if(in == 357) begin
					state<=2;
					out<=52;
				end
				if(in == 358) begin
					state<=2;
					out<=53;
				end
				if(in == 359) begin
					state<=2;
					out<=54;
				end
				if(in == 360) begin
					state<=2;
					out<=55;
				end
				if(in == 361) begin
					state<=2;
					out<=56;
				end
				if(in == 362) begin
					state<=2;
					out<=57;
				end
				if(in == 363) begin
					state<=2;
					out<=58;
				end
				if(in == 364) begin
					state<=2;
					out<=59;
				end
				if(in == 365) begin
					state<=2;
					out<=60;
				end
				if(in == 366) begin
					state<=2;
					out<=61;
				end
				if(in == 367) begin
					state<=2;
					out<=62;
				end
				if(in == 368) begin
					state<=2;
					out<=63;
				end
				if(in == 369) begin
					state<=2;
					out<=64;
				end
				if(in == 370) begin
					state<=2;
					out<=65;
				end
				if(in == 371) begin
					state<=2;
					out<=66;
				end
				if(in == 372) begin
					state<=2;
					out<=67;
				end
				if(in == 373) begin
					state<=2;
					out<=68;
				end
				if(in == 374) begin
					state<=2;
					out<=69;
				end
				if(in == 375) begin
					state<=2;
					out<=70;
				end
				if(in == 376) begin
					state<=2;
					out<=71;
				end
				if(in == 377) begin
					state<=2;
					out<=72;
				end
				if(in == 378) begin
					state<=2;
					out<=73;
				end
				if(in == 379) begin
					state<=2;
					out<=74;
				end
				if(in == 380) begin
					state<=2;
					out<=75;
				end
				if(in == 381) begin
					state<=2;
					out<=76;
				end
				if(in == 382) begin
					state<=2;
					out<=77;
				end
				if(in == 383) begin
					state<=2;
					out<=78;
				end
				if(in == 384) begin
					state<=2;
					out<=79;
				end
				if(in == 385) begin
					state<=2;
					out<=80;
				end
				if(in == 386) begin
					state<=2;
					out<=81;
				end
				if(in == 387) begin
					state<=2;
					out<=82;
				end
				if(in == 388) begin
					state<=2;
					out<=83;
				end
				if(in == 389) begin
					state<=2;
					out<=84;
				end
				if(in == 390) begin
					state<=2;
					out<=85;
				end
				if(in == 391) begin
					state<=2;
					out<=86;
				end
				if(in == 392) begin
					state<=2;
					out<=87;
				end
				if(in == 393) begin
					state<=2;
					out<=88;
				end
				if(in == 394) begin
					state<=2;
					out<=89;
				end
				if(in == 395) begin
					state<=2;
					out<=90;
				end
				if(in == 396) begin
					state<=2;
					out<=91;
				end
				if(in == 397) begin
					state<=2;
					out<=92;
				end
				if(in == 398) begin
					state<=2;
					out<=93;
				end
				if(in == 399) begin
					state<=2;
					out<=94;
				end
				if(in == 400) begin
					state<=2;
					out<=95;
				end
				if(in == 401) begin
					state<=2;
					out<=96;
				end
				if(in == 402) begin
					state<=2;
					out<=97;
				end
				if(in == 403) begin
					state<=2;
					out<=98;
				end
				if(in == 404) begin
					state<=2;
					out<=99;
				end
				if(in == 405) begin
					state<=2;
					out<=100;
				end
				if(in == 406) begin
					state<=2;
					out<=101;
				end
				if(in == 407) begin
					state<=2;
					out<=102;
				end
				if(in == 408) begin
					state<=2;
					out<=103;
				end
				if(in == 409) begin
					state<=2;
					out<=104;
				end
				if(in == 410) begin
					state<=2;
					out<=105;
				end
				if(in == 411) begin
					state<=2;
					out<=106;
				end
				if(in == 412) begin
					state<=2;
					out<=107;
				end
				if(in == 413) begin
					state<=2;
					out<=108;
				end
				if(in == 414) begin
					state<=2;
					out<=109;
				end
				if(in == 415) begin
					state<=2;
					out<=110;
				end
				if(in == 416) begin
					state<=2;
					out<=111;
				end
				if(in == 417) begin
					state<=2;
					out<=112;
				end
				if(in == 418) begin
					state<=2;
					out<=113;
				end
				if(in == 419) begin
					state<=2;
					out<=114;
				end
				if(in == 420) begin
					state<=2;
					out<=115;
				end
				if(in == 421) begin
					state<=2;
					out<=116;
				end
				if(in == 422) begin
					state<=2;
					out<=117;
				end
				if(in == 423) begin
					state<=2;
					out<=118;
				end
				if(in == 424) begin
					state<=2;
					out<=119;
				end
				if(in == 425) begin
					state<=2;
					out<=120;
				end
				if(in == 426) begin
					state<=2;
					out<=121;
				end
				if(in == 427) begin
					state<=2;
					out<=122;
				end
				if(in == 428) begin
					state<=2;
					out<=123;
				end
				if(in == 429) begin
					state<=2;
					out<=124;
				end
				if(in == 430) begin
					state<=2;
					out<=125;
				end
				if(in == 431) begin
					state<=2;
					out<=126;
				end
				if(in == 432) begin
					state<=2;
					out<=127;
				end
				if(in == 433) begin
					state<=2;
					out<=128;
				end
				if(in == 434) begin
					state<=2;
					out<=129;
				end
				if(in == 435) begin
					state<=2;
					out<=130;
				end
				if(in == 436) begin
					state<=2;
					out<=131;
				end
				if(in == 437) begin
					state<=2;
					out<=132;
				end
				if(in == 438) begin
					state<=2;
					out<=133;
				end
				if(in == 439) begin
					state<=2;
					out<=134;
				end
				if(in == 440) begin
					state<=2;
					out<=135;
				end
				if(in == 441) begin
					state<=2;
					out<=136;
				end
				if(in == 442) begin
					state<=2;
					out<=137;
				end
				if(in == 443) begin
					state<=2;
					out<=138;
				end
				if(in == 444) begin
					state<=2;
					out<=139;
				end
				if(in == 445) begin
					state<=2;
					out<=140;
				end
				if(in == 446) begin
					state<=2;
					out<=141;
				end
				if(in == 447) begin
					state<=2;
					out<=142;
				end
				if(in == 448) begin
					state<=2;
					out<=143;
				end
				if(in == 449) begin
					state<=2;
					out<=144;
				end
				if(in == 450) begin
					state<=2;
					out<=145;
				end
				if(in == 451) begin
					state<=2;
					out<=146;
				end
				if(in == 452) begin
					state<=2;
					out<=147;
				end
				if(in == 453) begin
					state<=2;
					out<=148;
				end
				if(in == 454) begin
					state<=2;
					out<=149;
				end
				if(in == 455) begin
					state<=2;
					out<=150;
				end
				if(in == 456) begin
					state<=2;
					out<=151;
				end
				if(in == 457) begin
					state<=2;
					out<=152;
				end
				if(in == 458) begin
					state<=2;
					out<=153;
				end
				if(in == 459) begin
					state<=2;
					out<=154;
				end
				if(in == 460) begin
					state<=2;
					out<=155;
				end
				if(in == 461) begin
					state<=2;
					out<=156;
				end
				if(in == 462) begin
					state<=2;
					out<=157;
				end
				if(in == 463) begin
					state<=2;
					out<=158;
				end
				if(in == 464) begin
					state<=2;
					out<=159;
				end
				if(in == 465) begin
					state<=2;
					out<=160;
				end
				if(in == 466) begin
					state<=2;
					out<=161;
				end
				if(in == 467) begin
					state<=2;
					out<=162;
				end
				if(in == 468) begin
					state<=2;
					out<=163;
				end
				if(in == 469) begin
					state<=2;
					out<=164;
				end
				if(in == 470) begin
					state<=2;
					out<=165;
				end
				if(in == 471) begin
					state<=2;
					out<=166;
				end
				if(in == 472) begin
					state<=2;
					out<=167;
				end
				if(in == 473) begin
					state<=2;
					out<=168;
				end
				if(in == 474) begin
					state<=2;
					out<=169;
				end
				if(in == 475) begin
					state<=2;
					out<=170;
				end
				if(in == 476) begin
					state<=2;
					out<=171;
				end
				if(in == 477) begin
					state<=2;
					out<=172;
				end
				if(in == 478) begin
					state<=2;
					out<=173;
				end
				if(in == 479) begin
					state<=2;
					out<=174;
				end
				if(in == 480) begin
					state<=2;
					out<=175;
				end
				if(in == 481) begin
					state<=2;
					out<=176;
				end
				if(in == 482) begin
					state<=2;
					out<=177;
				end
				if(in == 483) begin
					state<=2;
					out<=178;
				end
				if(in == 484) begin
					state<=2;
					out<=179;
				end
				if(in == 485) begin
					state<=2;
					out<=180;
				end
				if(in == 486) begin
					state<=2;
					out<=181;
				end
				if(in == 487) begin
					state<=2;
					out<=182;
				end
				if(in == 488) begin
					state<=2;
					out<=183;
				end
				if(in == 489) begin
					state<=2;
					out<=184;
				end
				if(in == 490) begin
					state<=2;
					out<=185;
				end
				if(in == 491) begin
					state<=2;
					out<=186;
				end
				if(in == 492) begin
					state<=2;
					out<=187;
				end
				if(in == 493) begin
					state<=2;
					out<=188;
				end
				if(in == 494) begin
					state<=2;
					out<=189;
				end
				if(in == 495) begin
					state<=2;
					out<=190;
				end
				if(in == 496) begin
					state<=2;
					out<=191;
				end
				if(in == 497) begin
					state<=2;
					out<=192;
				end
				if(in == 498) begin
					state<=2;
					out<=193;
				end
				if(in == 499) begin
					state<=2;
					out<=194;
				end
				if(in == 500) begin
					state<=2;
					out<=195;
				end
				if(in == 501) begin
					state<=2;
					out<=196;
				end
				if(in == 502) begin
					state<=2;
					out<=197;
				end
				if(in == 503) begin
					state<=2;
					out<=198;
				end
				if(in == 504) begin
					state<=2;
					out<=199;
				end
				if(in == 505) begin
					state<=2;
					out<=200;
				end
				if(in == 506) begin
					state<=2;
					out<=201;
				end
				if(in == 507) begin
					state<=2;
					out<=202;
				end
				if(in == 508) begin
					state<=2;
					out<=203;
				end
				if(in == 509) begin
					state<=2;
					out<=204;
				end
				if(in == 510) begin
					state<=2;
					out<=205;
				end
				if(in == 511) begin
					state<=2;
					out<=206;
				end
				if(in == 512) begin
					state<=2;
					out<=207;
				end
				if(in == 513) begin
					state<=2;
					out<=208;
				end
				if(in == 514) begin
					state<=2;
					out<=209;
				end
				if(in == 515) begin
					state<=2;
					out<=210;
				end
				if(in == 516) begin
					state<=2;
					out<=211;
				end
				if(in == 517) begin
					state<=2;
					out<=212;
				end
				if(in == 518) begin
					state<=2;
					out<=213;
				end
				if(in == 519) begin
					state<=2;
					out<=214;
				end
				if(in == 520) begin
					state<=2;
					out<=215;
				end
				if(in == 521) begin
					state<=2;
					out<=216;
				end
				if(in == 522) begin
					state<=2;
					out<=217;
				end
				if(in == 523) begin
					state<=2;
					out<=218;
				end
				if(in == 524) begin
					state<=2;
					out<=219;
				end
				if(in == 525) begin
					state<=2;
					out<=220;
				end
				if(in == 526) begin
					state<=2;
					out<=221;
				end
				if(in == 527) begin
					state<=2;
					out<=222;
				end
				if(in == 528) begin
					state<=2;
					out<=223;
				end
				if(in == 529) begin
					state<=2;
					out<=224;
				end
				if(in == 530) begin
					state<=2;
					out<=225;
				end
				if(in == 531) begin
					state<=2;
					out<=226;
				end
				if(in == 532) begin
					state<=2;
					out<=227;
				end
				if(in == 533) begin
					state<=2;
					out<=228;
				end
				if(in == 534) begin
					state<=2;
					out<=229;
				end
				if(in == 535) begin
					state<=2;
					out<=230;
				end
				if(in == 536) begin
					state<=2;
					out<=231;
				end
				if(in == 537) begin
					state<=2;
					out<=232;
				end
				if(in == 538) begin
					state<=2;
					out<=233;
				end
				if(in == 539) begin
					state<=2;
					out<=234;
				end
				if(in == 540) begin
					state<=2;
					out<=235;
				end
				if(in == 541) begin
					state<=2;
					out<=236;
				end
				if(in == 542) begin
					state<=2;
					out<=237;
				end
				if(in == 543) begin
					state<=2;
					out<=238;
				end
				if(in == 544) begin
					state<=2;
					out<=239;
				end
				if(in == 545) begin
					state<=2;
					out<=240;
				end
				if(in == 546) begin
					state<=2;
					out<=241;
				end
				if(in == 547) begin
					state<=2;
					out<=242;
				end
				if(in == 548) begin
					state<=2;
					out<=243;
				end
				if(in == 549) begin
					state<=2;
					out<=244;
				end
				if(in == 550) begin
					state<=2;
					out<=245;
				end
				if(in == 551) begin
					state<=2;
					out<=246;
				end
				if(in == 552) begin
					state<=2;
					out<=247;
				end
				if(in == 553) begin
					state<=2;
					out<=248;
				end
				if(in == 554) begin
					state<=2;
					out<=249;
				end
				if(in == 555) begin
					state<=2;
					out<=250;
				end
				if(in == 556) begin
					state<=2;
					out<=251;
				end
				if(in == 557) begin
					state<=2;
					out<=252;
				end
				if(in == 558) begin
					state<=2;
					out<=253;
				end
				if(in == 559) begin
					state<=2;
					out<=254;
				end
				if(in == 560) begin
					state<=2;
					out<=255;
				end
				if(in == 561) begin
					state<=2;
					out<=0;
				end
				if(in == 562) begin
					state<=2;
					out<=1;
				end
				if(in == 563) begin
					state<=2;
					out<=2;
				end
				if(in == 564) begin
					state<=2;
					out<=3;
				end
				if(in == 565) begin
					state<=2;
					out<=4;
				end
				if(in == 566) begin
					state<=2;
					out<=5;
				end
				if(in == 567) begin
					state<=2;
					out<=6;
				end
				if(in == 568) begin
					state<=2;
					out<=7;
				end
				if(in == 569) begin
					state<=2;
					out<=8;
				end
				if(in == 570) begin
					state<=2;
					out<=9;
				end
				if(in == 571) begin
					state<=2;
					out<=10;
				end
				if(in == 572) begin
					state<=2;
					out<=11;
				end
				if(in == 573) begin
					state<=2;
					out<=12;
				end
				if(in == 574) begin
					state<=2;
					out<=13;
				end
				if(in == 575) begin
					state<=2;
					out<=14;
				end
				if(in == 576) begin
					state<=2;
					out<=15;
				end
				if(in == 577) begin
					state<=2;
					out<=16;
				end
				if(in == 578) begin
					state<=2;
					out<=17;
				end
				if(in == 579) begin
					state<=2;
					out<=18;
				end
				if(in == 580) begin
					state<=2;
					out<=19;
				end
				if(in == 581) begin
					state<=2;
					out<=20;
				end
				if(in == 582) begin
					state<=2;
					out<=21;
				end
				if(in == 583) begin
					state<=2;
					out<=22;
				end
				if(in == 584) begin
					state<=2;
					out<=23;
				end
				if(in == 585) begin
					state<=2;
					out<=24;
				end
				if(in == 586) begin
					state<=2;
					out<=25;
				end
				if(in == 587) begin
					state<=2;
					out<=26;
				end
				if(in == 588) begin
					state<=2;
					out<=27;
				end
				if(in == 589) begin
					state<=2;
					out<=28;
				end
				if(in == 590) begin
					state<=2;
					out<=29;
				end
				if(in == 591) begin
					state<=2;
					out<=30;
				end
				if(in == 592) begin
					state<=2;
					out<=31;
				end
				if(in == 593) begin
					state<=2;
					out<=32;
				end
				if(in == 594) begin
					state<=2;
					out<=33;
				end
				if(in == 595) begin
					state<=2;
					out<=34;
				end
				if(in == 596) begin
					state<=2;
					out<=35;
				end
				if(in == 597) begin
					state<=2;
					out<=36;
				end
				if(in == 598) begin
					state<=2;
					out<=37;
				end
				if(in == 599) begin
					state<=2;
					out<=38;
				end
				if(in == 600) begin
					state<=2;
					out<=39;
				end
				if(in == 601) begin
					state<=2;
					out<=40;
				end
				if(in == 602) begin
					state<=2;
					out<=41;
				end
				if(in == 603) begin
					state<=2;
					out<=42;
				end
				if(in == 604) begin
					state<=2;
					out<=43;
				end
				if(in == 605) begin
					state<=2;
					out<=44;
				end
				if(in == 606) begin
					state<=2;
					out<=45;
				end
				if(in == 607) begin
					state<=2;
					out<=46;
				end
				if(in == 608) begin
					state<=2;
					out<=47;
				end
				if(in == 609) begin
					state<=2;
					out<=48;
				end
				if(in == 610) begin
					state<=2;
					out<=49;
				end
				if(in == 611) begin
					state<=2;
					out<=50;
				end
				if(in == 612) begin
					state<=2;
					out<=51;
				end
				if(in == 613) begin
					state<=2;
					out<=52;
				end
				if(in == 614) begin
					state<=2;
					out<=53;
				end
				if(in == 615) begin
					state<=2;
					out<=54;
				end
				if(in == 616) begin
					state<=2;
					out<=55;
				end
				if(in == 617) begin
					state<=2;
					out<=56;
				end
				if(in == 618) begin
					state<=2;
					out<=57;
				end
				if(in == 619) begin
					state<=2;
					out<=58;
				end
				if(in == 620) begin
					state<=2;
					out<=59;
				end
				if(in == 621) begin
					state<=2;
					out<=60;
				end
				if(in == 622) begin
					state<=2;
					out<=61;
				end
				if(in == 623) begin
					state<=2;
					out<=62;
				end
				if(in == 624) begin
					state<=2;
					out<=63;
				end
				if(in == 625) begin
					state<=2;
					out<=64;
				end
				if(in == 626) begin
					state<=2;
					out<=65;
				end
				if(in == 627) begin
					state<=2;
					out<=66;
				end
				if(in == 628) begin
					state<=2;
					out<=67;
				end
				if(in == 629) begin
					state<=2;
					out<=68;
				end
				if(in == 630) begin
					state<=2;
					out<=69;
				end
				if(in == 631) begin
					state<=2;
					out<=70;
				end
				if(in == 632) begin
					state<=2;
					out<=71;
				end
				if(in == 633) begin
					state<=2;
					out<=72;
				end
				if(in == 634) begin
					state<=2;
					out<=73;
				end
				if(in == 635) begin
					state<=2;
					out<=74;
				end
				if(in == 636) begin
					state<=2;
					out<=75;
				end
				if(in == 637) begin
					state<=2;
					out<=76;
				end
				if(in == 638) begin
					state<=2;
					out<=77;
				end
				if(in == 639) begin
					state<=2;
					out<=78;
				end
				if(in == 640) begin
					state<=2;
					out<=79;
				end
				if(in == 641) begin
					state<=2;
					out<=80;
				end
				if(in == 642) begin
					state<=2;
					out<=81;
				end
				if(in == 643) begin
					state<=2;
					out<=82;
				end
				if(in == 644) begin
					state<=2;
					out<=83;
				end
				if(in == 645) begin
					state<=2;
					out<=84;
				end
				if(in == 646) begin
					state<=2;
					out<=85;
				end
				if(in == 647) begin
					state<=2;
					out<=86;
				end
				if(in == 648) begin
					state<=2;
					out<=87;
				end
				if(in == 649) begin
					state<=2;
					out<=88;
				end
				if(in == 650) begin
					state<=2;
					out<=89;
				end
				if(in == 651) begin
					state<=2;
					out<=90;
				end
				if(in == 652) begin
					state<=2;
					out<=91;
				end
				if(in == 653) begin
					state<=2;
					out<=92;
				end
				if(in == 654) begin
					state<=2;
					out<=93;
				end
				if(in == 655) begin
					state<=2;
					out<=94;
				end
				if(in == 656) begin
					state<=2;
					out<=95;
				end
				if(in == 657) begin
					state<=2;
					out<=96;
				end
				if(in == 658) begin
					state<=2;
					out<=97;
				end
				if(in == 659) begin
					state<=2;
					out<=98;
				end
				if(in == 660) begin
					state<=2;
					out<=99;
				end
				if(in == 661) begin
					state<=2;
					out<=100;
				end
				if(in == 662) begin
					state<=2;
					out<=101;
				end
				if(in == 663) begin
					state<=2;
					out<=102;
				end
				if(in == 664) begin
					state<=2;
					out<=103;
				end
				if(in == 665) begin
					state<=2;
					out<=104;
				end
				if(in == 666) begin
					state<=2;
					out<=105;
				end
				if(in == 667) begin
					state<=2;
					out<=106;
				end
				if(in == 668) begin
					state<=2;
					out<=107;
				end
				if(in == 669) begin
					state<=2;
					out<=108;
				end
				if(in == 670) begin
					state<=2;
					out<=109;
				end
				if(in == 671) begin
					state<=2;
					out<=110;
				end
				if(in == 672) begin
					state<=2;
					out<=111;
				end
				if(in == 673) begin
					state<=2;
					out<=112;
				end
				if(in == 674) begin
					state<=2;
					out<=113;
				end
				if(in == 675) begin
					state<=2;
					out<=114;
				end
				if(in == 676) begin
					state<=2;
					out<=115;
				end
				if(in == 677) begin
					state<=2;
					out<=116;
				end
				if(in == 678) begin
					state<=2;
					out<=117;
				end
				if(in == 679) begin
					state<=2;
					out<=118;
				end
				if(in == 680) begin
					state<=2;
					out<=119;
				end
				if(in == 681) begin
					state<=2;
					out<=120;
				end
				if(in == 682) begin
					state<=2;
					out<=121;
				end
				if(in == 683) begin
					state<=2;
					out<=122;
				end
				if(in == 684) begin
					state<=2;
					out<=123;
				end
				if(in == 685) begin
					state<=2;
					out<=124;
				end
				if(in == 686) begin
					state<=2;
					out<=125;
				end
				if(in == 687) begin
					state<=2;
					out<=126;
				end
				if(in == 688) begin
					state<=2;
					out<=127;
				end
				if(in == 689) begin
					state<=2;
					out<=128;
				end
				if(in == 690) begin
					state<=2;
					out<=129;
				end
				if(in == 691) begin
					state<=2;
					out<=130;
				end
				if(in == 692) begin
					state<=2;
					out<=131;
				end
				if(in == 693) begin
					state<=2;
					out<=132;
				end
				if(in == 694) begin
					state<=2;
					out<=133;
				end
				if(in == 695) begin
					state<=2;
					out<=134;
				end
				if(in == 696) begin
					state<=2;
					out<=135;
				end
				if(in == 697) begin
					state<=2;
					out<=136;
				end
				if(in == 698) begin
					state<=2;
					out<=137;
				end
				if(in == 699) begin
					state<=2;
					out<=138;
				end
				if(in == 700) begin
					state<=2;
					out<=139;
				end
				if(in == 701) begin
					state<=2;
					out<=140;
				end
				if(in == 702) begin
					state<=2;
					out<=141;
				end
				if(in == 703) begin
					state<=2;
					out<=142;
				end
				if(in == 704) begin
					state<=2;
					out<=143;
				end
				if(in == 705) begin
					state<=2;
					out<=144;
				end
				if(in == 706) begin
					state<=2;
					out<=145;
				end
				if(in == 707) begin
					state<=2;
					out<=146;
				end
				if(in == 708) begin
					state<=2;
					out<=147;
				end
				if(in == 709) begin
					state<=2;
					out<=148;
				end
				if(in == 710) begin
					state<=2;
					out<=149;
				end
				if(in == 711) begin
					state<=2;
					out<=150;
				end
				if(in == 712) begin
					state<=2;
					out<=151;
				end
				if(in == 713) begin
					state<=2;
					out<=152;
				end
				if(in == 714) begin
					state<=2;
					out<=153;
				end
				if(in == 715) begin
					state<=2;
					out<=154;
				end
				if(in == 716) begin
					state<=2;
					out<=155;
				end
				if(in == 717) begin
					state<=2;
					out<=156;
				end
				if(in == 718) begin
					state<=2;
					out<=157;
				end
				if(in == 719) begin
					state<=2;
					out<=158;
				end
				if(in == 720) begin
					state<=2;
					out<=159;
				end
				if(in == 721) begin
					state<=2;
					out<=160;
				end
				if(in == 722) begin
					state<=2;
					out<=161;
				end
				if(in == 723) begin
					state<=2;
					out<=162;
				end
				if(in == 724) begin
					state<=2;
					out<=163;
				end
				if(in == 725) begin
					state<=2;
					out<=164;
				end
				if(in == 726) begin
					state<=2;
					out<=165;
				end
				if(in == 727) begin
					state<=2;
					out<=166;
				end
				if(in == 728) begin
					state<=2;
					out<=167;
				end
				if(in == 729) begin
					state<=2;
					out<=168;
				end
				if(in == 730) begin
					state<=2;
					out<=169;
				end
				if(in == 731) begin
					state<=2;
					out<=170;
				end
				if(in == 732) begin
					state<=2;
					out<=171;
				end
				if(in == 733) begin
					state<=2;
					out<=172;
				end
				if(in == 734) begin
					state<=2;
					out<=173;
				end
				if(in == 735) begin
					state<=2;
					out<=174;
				end
				if(in == 736) begin
					state<=2;
					out<=175;
				end
				if(in == 737) begin
					state<=2;
					out<=176;
				end
				if(in == 738) begin
					state<=2;
					out<=177;
				end
				if(in == 739) begin
					state<=2;
					out<=178;
				end
				if(in == 740) begin
					state<=2;
					out<=179;
				end
				if(in == 741) begin
					state<=2;
					out<=180;
				end
				if(in == 742) begin
					state<=2;
					out<=181;
				end
				if(in == 743) begin
					state<=2;
					out<=182;
				end
				if(in == 744) begin
					state<=2;
					out<=183;
				end
				if(in == 745) begin
					state<=2;
					out<=184;
				end
				if(in == 746) begin
					state<=2;
					out<=185;
				end
				if(in == 747) begin
					state<=2;
					out<=186;
				end
				if(in == 748) begin
					state<=2;
					out<=187;
				end
				if(in == 749) begin
					state<=2;
					out<=188;
				end
				if(in == 750) begin
					state<=2;
					out<=189;
				end
				if(in == 751) begin
					state<=2;
					out<=190;
				end
				if(in == 752) begin
					state<=2;
					out<=191;
				end
				if(in == 753) begin
					state<=2;
					out<=192;
				end
				if(in == 754) begin
					state<=2;
					out<=193;
				end
				if(in == 755) begin
					state<=2;
					out<=194;
				end
				if(in == 756) begin
					state<=2;
					out<=195;
				end
				if(in == 757) begin
					state<=2;
					out<=196;
				end
				if(in == 758) begin
					state<=2;
					out<=197;
				end
				if(in == 759) begin
					state<=2;
					out<=198;
				end
				if(in == 760) begin
					state<=2;
					out<=199;
				end
				if(in == 761) begin
					state<=2;
					out<=200;
				end
				if(in == 762) begin
					state<=2;
					out<=201;
				end
				if(in == 763) begin
					state<=2;
					out<=202;
				end
				if(in == 764) begin
					state<=2;
					out<=203;
				end
				if(in == 765) begin
					state<=2;
					out<=204;
				end
				if(in == 766) begin
					state<=2;
					out<=205;
				end
				if(in == 767) begin
					state<=2;
					out<=206;
				end
				if(in == 768) begin
					state<=2;
					out<=207;
				end
				if(in == 769) begin
					state<=2;
					out<=208;
				end
				if(in == 770) begin
					state<=2;
					out<=209;
				end
				if(in == 771) begin
					state<=2;
					out<=210;
				end
				if(in == 772) begin
					state<=2;
					out<=211;
				end
				if(in == 773) begin
					state<=2;
					out<=212;
				end
				if(in == 774) begin
					state<=2;
					out<=213;
				end
				if(in == 775) begin
					state<=2;
					out<=214;
				end
				if(in == 776) begin
					state<=2;
					out<=215;
				end
				if(in == 777) begin
					state<=2;
					out<=216;
				end
				if(in == 778) begin
					state<=2;
					out<=217;
				end
				if(in == 779) begin
					state<=2;
					out<=218;
				end
				if(in == 780) begin
					state<=2;
					out<=219;
				end
				if(in == 781) begin
					state<=2;
					out<=220;
				end
				if(in == 782) begin
					state<=2;
					out<=221;
				end
				if(in == 783) begin
					state<=2;
					out<=222;
				end
				if(in == 784) begin
					state<=2;
					out<=223;
				end
				if(in == 785) begin
					state<=2;
					out<=224;
				end
				if(in == 786) begin
					state<=2;
					out<=225;
				end
				if(in == 787) begin
					state<=2;
					out<=226;
				end
				if(in == 788) begin
					state<=2;
					out<=227;
				end
				if(in == 789) begin
					state<=2;
					out<=228;
				end
				if(in == 790) begin
					state<=2;
					out<=229;
				end
				if(in == 791) begin
					state<=2;
					out<=230;
				end
				if(in == 792) begin
					state<=2;
					out<=231;
				end
				if(in == 793) begin
					state<=2;
					out<=232;
				end
				if(in == 794) begin
					state<=2;
					out<=233;
				end
				if(in == 795) begin
					state<=2;
					out<=234;
				end
				if(in == 796) begin
					state<=2;
					out<=235;
				end
				if(in == 797) begin
					state<=2;
					out<=236;
				end
				if(in == 798) begin
					state<=2;
					out<=237;
				end
				if(in == 799) begin
					state<=2;
					out<=238;
				end
				if(in == 800) begin
					state<=2;
					out<=239;
				end
				if(in == 801) begin
					state<=2;
					out<=240;
				end
				if(in == 802) begin
					state<=2;
					out<=241;
				end
				if(in == 803) begin
					state<=2;
					out<=242;
				end
				if(in == 804) begin
					state<=2;
					out<=243;
				end
				if(in == 805) begin
					state<=2;
					out<=244;
				end
				if(in == 806) begin
					state<=2;
					out<=245;
				end
				if(in == 807) begin
					state<=2;
					out<=246;
				end
				if(in == 808) begin
					state<=2;
					out<=247;
				end
				if(in == 809) begin
					state<=2;
					out<=248;
				end
				if(in == 810) begin
					state<=2;
					out<=249;
				end
				if(in == 811) begin
					state<=2;
					out<=250;
				end
				if(in == 812) begin
					state<=2;
					out<=251;
				end
				if(in == 813) begin
					state<=2;
					out<=252;
				end
				if(in == 814) begin
					state<=2;
					out<=253;
				end
				if(in == 815) begin
					state<=2;
					out<=254;
				end
				if(in == 816) begin
					state<=2;
					out<=255;
				end
				if(in == 817) begin
					state<=2;
					out<=0;
				end
				if(in == 818) begin
					state<=2;
					out<=1;
				end
				if(in == 819) begin
					state<=2;
					out<=2;
				end
				if(in == 820) begin
					state<=2;
					out<=3;
				end
				if(in == 821) begin
					state<=2;
					out<=4;
				end
				if(in == 822) begin
					state<=2;
					out<=5;
				end
				if(in == 823) begin
					state<=2;
					out<=6;
				end
				if(in == 824) begin
					state<=2;
					out<=7;
				end
				if(in == 825) begin
					state<=2;
					out<=8;
				end
				if(in == 826) begin
					state<=2;
					out<=9;
				end
				if(in == 827) begin
					state<=2;
					out<=10;
				end
				if(in == 828) begin
					state<=2;
					out<=11;
				end
				if(in == 829) begin
					state<=2;
					out<=12;
				end
				if(in == 830) begin
					state<=2;
					out<=13;
				end
				if(in == 831) begin
					state<=2;
					out<=14;
				end
				if(in == 832) begin
					state<=2;
					out<=15;
				end
				if(in == 833) begin
					state<=2;
					out<=16;
				end
				if(in == 834) begin
					state<=2;
					out<=17;
				end
				if(in == 835) begin
					state<=2;
					out<=18;
				end
				if(in == 836) begin
					state<=2;
					out<=19;
				end
				if(in == 837) begin
					state<=2;
					out<=20;
				end
				if(in == 838) begin
					state<=2;
					out<=21;
				end
				if(in == 839) begin
					state<=2;
					out<=22;
				end
				if(in == 840) begin
					state<=2;
					out<=23;
				end
				if(in == 841) begin
					state<=2;
					out<=24;
				end
				if(in == 842) begin
					state<=2;
					out<=25;
				end
				if(in == 843) begin
					state<=2;
					out<=26;
				end
				if(in == 844) begin
					state<=2;
					out<=27;
				end
				if(in == 845) begin
					state<=2;
					out<=28;
				end
				if(in == 846) begin
					state<=2;
					out<=29;
				end
				if(in == 847) begin
					state<=2;
					out<=30;
				end
				if(in == 848) begin
					state<=2;
					out<=31;
				end
				if(in == 849) begin
					state<=2;
					out<=32;
				end
				if(in == 850) begin
					state<=2;
					out<=33;
				end
				if(in == 851) begin
					state<=2;
					out<=34;
				end
				if(in == 852) begin
					state<=2;
					out<=35;
				end
				if(in == 853) begin
					state<=2;
					out<=36;
				end
				if(in == 854) begin
					state<=2;
					out<=37;
				end
				if(in == 855) begin
					state<=2;
					out<=38;
				end
				if(in == 856) begin
					state<=2;
					out<=39;
				end
				if(in == 857) begin
					state<=2;
					out<=40;
				end
				if(in == 858) begin
					state<=2;
					out<=41;
				end
				if(in == 859) begin
					state<=2;
					out<=42;
				end
				if(in == 860) begin
					state<=2;
					out<=43;
				end
				if(in == 861) begin
					state<=2;
					out<=44;
				end
				if(in == 862) begin
					state<=2;
					out<=45;
				end
				if(in == 863) begin
					state<=2;
					out<=46;
				end
				if(in == 864) begin
					state<=2;
					out<=47;
				end
				if(in == 865) begin
					state<=2;
					out<=48;
				end
				if(in == 866) begin
					state<=2;
					out<=49;
				end
				if(in == 867) begin
					state<=2;
					out<=50;
				end
				if(in == 868) begin
					state<=2;
					out<=51;
				end
				if(in == 869) begin
					state<=2;
					out<=52;
				end
				if(in == 870) begin
					state<=2;
					out<=53;
				end
				if(in == 871) begin
					state<=2;
					out<=54;
				end
				if(in == 872) begin
					state<=2;
					out<=55;
				end
				if(in == 873) begin
					state<=2;
					out<=56;
				end
				if(in == 874) begin
					state<=2;
					out<=57;
				end
				if(in == 875) begin
					state<=2;
					out<=58;
				end
				if(in == 876) begin
					state<=2;
					out<=59;
				end
				if(in == 877) begin
					state<=2;
					out<=60;
				end
				if(in == 878) begin
					state<=2;
					out<=61;
				end
				if(in == 879) begin
					state<=2;
					out<=62;
				end
				if(in == 880) begin
					state<=2;
					out<=63;
				end
				if(in == 881) begin
					state<=2;
					out<=64;
				end
				if(in == 882) begin
					state<=2;
					out<=65;
				end
				if(in == 883) begin
					state<=2;
					out<=66;
				end
				if(in == 884) begin
					state<=2;
					out<=67;
				end
				if(in == 885) begin
					state<=2;
					out<=68;
				end
				if(in == 886) begin
					state<=2;
					out<=69;
				end
				if(in == 887) begin
					state<=2;
					out<=70;
				end
				if(in == 888) begin
					state<=2;
					out<=71;
				end
				if(in == 889) begin
					state<=2;
					out<=72;
				end
				if(in == 890) begin
					state<=2;
					out<=73;
				end
				if(in == 891) begin
					state<=2;
					out<=74;
				end
				if(in == 892) begin
					state<=2;
					out<=75;
				end
				if(in == 893) begin
					state<=2;
					out<=76;
				end
				if(in == 894) begin
					state<=2;
					out<=77;
				end
				if(in == 895) begin
					state<=2;
					out<=78;
				end
				if(in == 896) begin
					state<=2;
					out<=79;
				end
				if(in == 897) begin
					state<=2;
					out<=80;
				end
				if(in == 898) begin
					state<=2;
					out<=81;
				end
				if(in == 899) begin
					state<=2;
					out<=82;
				end
				if(in == 900) begin
					state<=2;
					out<=83;
				end
				if(in == 901) begin
					state<=2;
					out<=84;
				end
				if(in == 902) begin
					state<=2;
					out<=85;
				end
				if(in == 903) begin
					state<=2;
					out<=86;
				end
				if(in == 904) begin
					state<=2;
					out<=87;
				end
				if(in == 905) begin
					state<=2;
					out<=88;
				end
				if(in == 906) begin
					state<=2;
					out<=89;
				end
				if(in == 907) begin
					state<=2;
					out<=90;
				end
				if(in == 908) begin
					state<=2;
					out<=91;
				end
				if(in == 909) begin
					state<=2;
					out<=92;
				end
				if(in == 910) begin
					state<=2;
					out<=93;
				end
				if(in == 911) begin
					state<=2;
					out<=94;
				end
				if(in == 912) begin
					state<=2;
					out<=95;
				end
				if(in == 913) begin
					state<=2;
					out<=96;
				end
				if(in == 914) begin
					state<=2;
					out<=97;
				end
				if(in == 915) begin
					state<=2;
					out<=98;
				end
				if(in == 916) begin
					state<=2;
					out<=99;
				end
				if(in == 917) begin
					state<=2;
					out<=100;
				end
				if(in == 918) begin
					state<=2;
					out<=101;
				end
				if(in == 919) begin
					state<=2;
					out<=102;
				end
				if(in == 920) begin
					state<=2;
					out<=103;
				end
				if(in == 921) begin
					state<=2;
					out<=104;
				end
				if(in == 922) begin
					state<=2;
					out<=105;
				end
				if(in == 923) begin
					state<=2;
					out<=106;
				end
				if(in == 924) begin
					state<=2;
					out<=107;
				end
				if(in == 925) begin
					state<=2;
					out<=108;
				end
				if(in == 926) begin
					state<=2;
					out<=109;
				end
				if(in == 927) begin
					state<=2;
					out<=110;
				end
				if(in == 928) begin
					state<=2;
					out<=111;
				end
			end
			16: begin
				if(in == 0) begin
					state<=16;
					out<=112;
				end
				if(in == 1) begin
					state<=1;
					out<=113;
				end
				if(in == 2) begin
					state<=16;
					out<=114;
				end
				if(in == 3) begin
					state<=16;
					out<=115;
				end
				if(in == 4) begin
					state<=16;
					out<=116;
				end
				if(in == 5) begin
					state<=16;
					out<=117;
				end
				if(in == 6) begin
					state<=16;
					out<=118;
				end
				if(in == 7) begin
					state<=16;
					out<=119;
				end
				if(in == 8) begin
					state<=16;
					out<=120;
				end
				if(in == 9) begin
					state<=16;
					out<=121;
				end
				if(in == 10) begin
					state<=16;
					out<=122;
				end
				if(in == 11) begin
					state<=16;
					out<=123;
				end
				if(in == 12) begin
					state<=16;
					out<=124;
				end
				if(in == 13) begin
					state<=16;
					out<=125;
				end
				if(in == 14) begin
					state<=16;
					out<=126;
				end
				if(in == 15) begin
					state<=16;
					out<=127;
				end
				if(in == 16) begin
					state<=16;
					out<=128;
				end
				if(in == 17) begin
					state<=16;
					out<=129;
				end
				if(in == 18) begin
					state<=16;
					out<=130;
				end
				if(in == 19) begin
					state<=16;
					out<=131;
				end
				if(in == 20) begin
					state<=16;
					out<=132;
				end
				if(in == 21) begin
					state<=16;
					out<=133;
				end
				if(in == 22) begin
					state<=16;
					out<=134;
				end
				if(in == 23) begin
					state<=16;
					out<=135;
				end
				if(in == 24) begin
					state<=16;
					out<=136;
				end
				if(in == 25) begin
					state<=16;
					out<=137;
				end
				if(in == 26) begin
					state<=16;
					out<=138;
				end
				if(in == 27) begin
					state<=16;
					out<=139;
				end
				if(in == 28) begin
					state<=16;
					out<=140;
				end
				if(in == 29) begin
					state<=16;
					out<=141;
				end
				if(in == 30) begin
					state<=16;
					out<=142;
				end
				if(in == 31) begin
					state<=16;
					out<=143;
				end
				if(in == 32) begin
					state<=16;
					out<=144;
				end
				if(in == 33) begin
					state<=16;
					out<=145;
				end
				if(in == 34) begin
					state<=16;
					out<=146;
				end
				if(in == 35) begin
					state<=16;
					out<=147;
				end
				if(in == 36) begin
					state<=16;
					out<=148;
				end
				if(in == 37) begin
					state<=16;
					out<=149;
				end
				if(in == 38) begin
					state<=16;
					out<=150;
				end
				if(in == 39) begin
					state<=16;
					out<=151;
				end
				if(in == 40) begin
					state<=16;
					out<=152;
				end
				if(in == 41) begin
					state<=16;
					out<=153;
				end
				if(in == 42) begin
					state<=16;
					out<=154;
				end
				if(in == 43) begin
					state<=16;
					out<=155;
				end
				if(in == 44) begin
					state<=16;
					out<=156;
				end
				if(in == 45) begin
					state<=16;
					out<=157;
				end
				if(in == 46) begin
					state<=16;
					out<=158;
				end
				if(in == 47) begin
					state<=16;
					out<=159;
				end
				if(in == 48) begin
					state<=16;
					out<=160;
				end
				if(in == 49) begin
					state<=16;
					out<=161;
				end
				if(in == 50) begin
					state<=16;
					out<=162;
				end
				if(in == 51) begin
					state<=16;
					out<=163;
				end
				if(in == 52) begin
					state<=16;
					out<=164;
				end
				if(in == 53) begin
					state<=16;
					out<=165;
				end
				if(in == 54) begin
					state<=16;
					out<=166;
				end
				if(in == 55) begin
					state<=16;
					out<=167;
				end
				if(in == 56) begin
					state<=16;
					out<=168;
				end
				if(in == 57) begin
					state<=16;
					out<=169;
				end
				if(in == 58) begin
					state<=16;
					out<=170;
				end
				if(in == 59) begin
					state<=16;
					out<=171;
				end
				if(in == 60) begin
					state<=16;
					out<=172;
				end
				if(in == 61) begin
					state<=16;
					out<=173;
				end
				if(in == 62) begin
					state<=16;
					out<=174;
				end
				if(in == 63) begin
					state<=16;
					out<=175;
				end
				if(in == 64) begin
					state<=16;
					out<=176;
				end
				if(in == 65) begin
					state<=16;
					out<=177;
				end
				if(in == 66) begin
					state<=16;
					out<=178;
				end
				if(in == 67) begin
					state<=16;
					out<=179;
				end
				if(in == 68) begin
					state<=16;
					out<=180;
				end
				if(in == 69) begin
					state<=16;
					out<=181;
				end
				if(in == 70) begin
					state<=16;
					out<=182;
				end
				if(in == 71) begin
					state<=16;
					out<=183;
				end
				if(in == 72) begin
					state<=16;
					out<=184;
				end
				if(in == 73) begin
					state<=16;
					out<=185;
				end
				if(in == 74) begin
					state<=16;
					out<=186;
				end
				if(in == 75) begin
					state<=16;
					out<=187;
				end
				if(in == 76) begin
					state<=16;
					out<=188;
				end
				if(in == 77) begin
					state<=16;
					out<=189;
				end
				if(in == 78) begin
					state<=16;
					out<=190;
				end
				if(in == 79) begin
					state<=16;
					out<=191;
				end
				if(in == 80) begin
					state<=16;
					out<=192;
				end
				if(in == 81) begin
					state<=16;
					out<=193;
				end
				if(in == 82) begin
					state<=16;
					out<=194;
				end
				if(in == 83) begin
					state<=16;
					out<=195;
				end
				if(in == 84) begin
					state<=16;
					out<=196;
				end
				if(in == 85) begin
					state<=16;
					out<=197;
				end
				if(in == 86) begin
					state<=16;
					out<=198;
				end
				if(in == 87) begin
					state<=16;
					out<=199;
				end
				if(in == 88) begin
					state<=16;
					out<=200;
				end
				if(in == 89) begin
					state<=16;
					out<=201;
				end
				if(in == 90) begin
					state<=16;
					out<=202;
				end
				if(in == 91) begin
					state<=16;
					out<=203;
				end
				if(in == 92) begin
					state<=16;
					out<=204;
				end
				if(in == 93) begin
					state<=16;
					out<=205;
				end
				if(in == 94) begin
					state<=16;
					out<=206;
				end
				if(in == 95) begin
					state<=16;
					out<=207;
				end
				if(in == 96) begin
					state<=16;
					out<=208;
				end
				if(in == 97) begin
					state<=16;
					out<=209;
				end
				if(in == 98) begin
					state<=16;
					out<=210;
				end
				if(in == 99) begin
					state<=16;
					out<=211;
				end
				if(in == 100) begin
					state<=16;
					out<=212;
				end
				if(in == 101) begin
					state<=16;
					out<=213;
				end
				if(in == 102) begin
					state<=16;
					out<=214;
				end
				if(in == 103) begin
					state<=16;
					out<=215;
				end
				if(in == 104) begin
					state<=16;
					out<=216;
				end
				if(in == 105) begin
					state<=16;
					out<=217;
				end
				if(in == 106) begin
					state<=16;
					out<=218;
				end
				if(in == 107) begin
					state<=16;
					out<=219;
				end
				if(in == 108) begin
					state<=16;
					out<=220;
				end
				if(in == 109) begin
					state<=16;
					out<=221;
				end
				if(in == 110) begin
					state<=16;
					out<=222;
				end
				if(in == 111) begin
					state<=16;
					out<=223;
				end
				if(in == 112) begin
					state<=16;
					out<=224;
				end
				if(in == 113) begin
					state<=16;
					out<=225;
				end
				if(in == 114) begin
					state<=16;
					out<=226;
				end
				if(in == 115) begin
					state<=16;
					out<=227;
				end
				if(in == 116) begin
					state<=16;
					out<=228;
				end
				if(in == 117) begin
					state<=16;
					out<=229;
				end
				if(in == 118) begin
					state<=16;
					out<=230;
				end
				if(in == 119) begin
					state<=16;
					out<=231;
				end
				if(in == 120) begin
					state<=16;
					out<=232;
				end
				if(in == 121) begin
					state<=16;
					out<=233;
				end
				if(in == 122) begin
					state<=16;
					out<=234;
				end
				if(in == 123) begin
					state<=16;
					out<=235;
				end
				if(in == 124) begin
					state<=16;
					out<=236;
				end
				if(in == 125) begin
					state<=16;
					out<=237;
				end
				if(in == 126) begin
					state<=16;
					out<=238;
				end
				if(in == 127) begin
					state<=16;
					out<=239;
				end
				if(in == 128) begin
					state<=16;
					out<=240;
				end
				if(in == 129) begin
					state<=16;
					out<=241;
				end
				if(in == 130) begin
					state<=16;
					out<=242;
				end
				if(in == 131) begin
					state<=16;
					out<=243;
				end
				if(in == 132) begin
					state<=16;
					out<=244;
				end
				if(in == 133) begin
					state<=16;
					out<=245;
				end
				if(in == 134) begin
					state<=16;
					out<=246;
				end
				if(in == 135) begin
					state<=16;
					out<=247;
				end
				if(in == 136) begin
					state<=16;
					out<=248;
				end
				if(in == 137) begin
					state<=16;
					out<=249;
				end
				if(in == 138) begin
					state<=16;
					out<=250;
				end
				if(in == 139) begin
					state<=16;
					out<=251;
				end
				if(in == 140) begin
					state<=16;
					out<=252;
				end
				if(in == 141) begin
					state<=16;
					out<=253;
				end
				if(in == 142) begin
					state<=16;
					out<=254;
				end
				if(in == 143) begin
					state<=16;
					out<=255;
				end
				if(in == 144) begin
					state<=16;
					out<=0;
				end
				if(in == 145) begin
					state<=16;
					out<=1;
				end
				if(in == 146) begin
					state<=16;
					out<=2;
				end
				if(in == 147) begin
					state<=16;
					out<=3;
				end
				if(in == 148) begin
					state<=16;
					out<=4;
				end
				if(in == 149) begin
					state<=16;
					out<=5;
				end
				if(in == 150) begin
					state<=16;
					out<=6;
				end
				if(in == 151) begin
					state<=16;
					out<=7;
				end
				if(in == 152) begin
					state<=16;
					out<=8;
				end
				if(in == 153) begin
					state<=16;
					out<=9;
				end
				if(in == 154) begin
					state<=16;
					out<=10;
				end
				if(in == 155) begin
					state<=16;
					out<=11;
				end
				if(in == 156) begin
					state<=16;
					out<=12;
				end
				if(in == 157) begin
					state<=16;
					out<=13;
				end
				if(in == 158) begin
					state<=16;
					out<=14;
				end
				if(in == 159) begin
					state<=16;
					out<=15;
				end
				if(in == 160) begin
					state<=16;
					out<=16;
				end
				if(in == 161) begin
					state<=16;
					out<=17;
				end
				if(in == 162) begin
					state<=16;
					out<=18;
				end
				if(in == 163) begin
					state<=16;
					out<=19;
				end
				if(in == 164) begin
					state<=16;
					out<=20;
				end
				if(in == 165) begin
					state<=16;
					out<=21;
				end
				if(in == 166) begin
					state<=16;
					out<=22;
				end
				if(in == 167) begin
					state<=16;
					out<=23;
				end
				if(in == 168) begin
					state<=16;
					out<=24;
				end
				if(in == 169) begin
					state<=16;
					out<=25;
				end
				if(in == 170) begin
					state<=16;
					out<=26;
				end
				if(in == 171) begin
					state<=16;
					out<=27;
				end
				if(in == 172) begin
					state<=16;
					out<=28;
				end
				if(in == 173) begin
					state<=16;
					out<=29;
				end
				if(in == 174) begin
					state<=16;
					out<=30;
				end
				if(in == 175) begin
					state<=16;
					out<=31;
				end
				if(in == 176) begin
					state<=16;
					out<=32;
				end
				if(in == 177) begin
					state<=16;
					out<=33;
				end
				if(in == 178) begin
					state<=16;
					out<=34;
				end
				if(in == 179) begin
					state<=16;
					out<=35;
				end
				if(in == 180) begin
					state<=16;
					out<=36;
				end
				if(in == 181) begin
					state<=16;
					out<=37;
				end
				if(in == 182) begin
					state<=16;
					out<=38;
				end
				if(in == 183) begin
					state<=16;
					out<=39;
				end
				if(in == 184) begin
					state<=16;
					out<=40;
				end
				if(in == 185) begin
					state<=16;
					out<=41;
				end
				if(in == 186) begin
					state<=16;
					out<=42;
				end
				if(in == 187) begin
					state<=16;
					out<=43;
				end
				if(in == 188) begin
					state<=16;
					out<=44;
				end
				if(in == 189) begin
					state<=16;
					out<=45;
				end
				if(in == 190) begin
					state<=16;
					out<=46;
				end
				if(in == 191) begin
					state<=16;
					out<=47;
				end
				if(in == 192) begin
					state<=16;
					out<=48;
				end
				if(in == 193) begin
					state<=16;
					out<=49;
				end
				if(in == 194) begin
					state<=16;
					out<=50;
				end
				if(in == 195) begin
					state<=16;
					out<=51;
				end
				if(in == 196) begin
					state<=16;
					out<=52;
				end
				if(in == 197) begin
					state<=16;
					out<=53;
				end
				if(in == 198) begin
					state<=16;
					out<=54;
				end
				if(in == 199) begin
					state<=16;
					out<=55;
				end
				if(in == 200) begin
					state<=16;
					out<=56;
				end
				if(in == 201) begin
					state<=16;
					out<=57;
				end
				if(in == 202) begin
					state<=16;
					out<=58;
				end
				if(in == 203) begin
					state<=16;
					out<=59;
				end
				if(in == 204) begin
					state<=16;
					out<=60;
				end
				if(in == 205) begin
					state<=16;
					out<=61;
				end
				if(in == 206) begin
					state<=16;
					out<=62;
				end
				if(in == 207) begin
					state<=16;
					out<=63;
				end
				if(in == 208) begin
					state<=16;
					out<=64;
				end
				if(in == 209) begin
					state<=16;
					out<=65;
				end
				if(in == 210) begin
					state<=16;
					out<=66;
				end
				if(in == 211) begin
					state<=16;
					out<=67;
				end
				if(in == 212) begin
					state<=16;
					out<=68;
				end
				if(in == 213) begin
					state<=16;
					out<=69;
				end
				if(in == 214) begin
					state<=16;
					out<=70;
				end
				if(in == 215) begin
					state<=16;
					out<=71;
				end
				if(in == 216) begin
					state<=16;
					out<=72;
				end
				if(in == 217) begin
					state<=16;
					out<=73;
				end
				if(in == 218) begin
					state<=16;
					out<=74;
				end
				if(in == 219) begin
					state<=16;
					out<=75;
				end
				if(in == 220) begin
					state<=16;
					out<=76;
				end
				if(in == 221) begin
					state<=16;
					out<=77;
				end
				if(in == 222) begin
					state<=16;
					out<=78;
				end
				if(in == 223) begin
					state<=16;
					out<=79;
				end
				if(in == 224) begin
					state<=16;
					out<=80;
				end
				if(in == 225) begin
					state<=16;
					out<=81;
				end
				if(in == 226) begin
					state<=16;
					out<=82;
				end
				if(in == 227) begin
					state<=16;
					out<=83;
				end
				if(in == 228) begin
					state<=16;
					out<=84;
				end
				if(in == 229) begin
					state<=16;
					out<=85;
				end
				if(in == 230) begin
					state<=16;
					out<=86;
				end
				if(in == 231) begin
					state<=16;
					out<=87;
				end
				if(in == 232) begin
					state<=16;
					out<=88;
				end
				if(in == 233) begin
					state<=16;
					out<=89;
				end
				if(in == 234) begin
					state<=16;
					out<=90;
				end
				if(in == 235) begin
					state<=16;
					out<=91;
				end
				if(in == 236) begin
					state<=16;
					out<=92;
				end
				if(in == 237) begin
					state<=16;
					out<=93;
				end
				if(in == 238) begin
					state<=16;
					out<=94;
				end
				if(in == 239) begin
					state<=16;
					out<=95;
				end
				if(in == 240) begin
					state<=16;
					out<=96;
				end
				if(in == 241) begin
					state<=16;
					out<=97;
				end
				if(in == 242) begin
					state<=16;
					out<=98;
				end
				if(in == 243) begin
					state<=16;
					out<=99;
				end
				if(in == 244) begin
					state<=16;
					out<=100;
				end
				if(in == 245) begin
					state<=16;
					out<=101;
				end
				if(in == 246) begin
					state<=16;
					out<=102;
				end
				if(in == 247) begin
					state<=16;
					out<=103;
				end
				if(in == 248) begin
					state<=16;
					out<=104;
				end
				if(in == 249) begin
					state<=16;
					out<=105;
				end
				if(in == 250) begin
					state<=16;
					out<=106;
				end
				if(in == 251) begin
					state<=16;
					out<=107;
				end
				if(in == 252) begin
					state<=16;
					out<=108;
				end
				if(in == 253) begin
					state<=16;
					out<=109;
				end
				if(in == 254) begin
					state<=16;
					out<=110;
				end
				if(in == 255) begin
					state<=16;
					out<=111;
				end
				if(in == 256) begin
					state<=16;
					out<=112;
				end
				if(in == 257) begin
					state<=16;
					out<=113;
				end
				if(in == 258) begin
					state<=16;
					out<=114;
				end
				if(in == 259) begin
					state<=16;
					out<=115;
				end
				if(in == 260) begin
					state<=16;
					out<=116;
				end
				if(in == 261) begin
					state<=16;
					out<=117;
				end
				if(in == 262) begin
					state<=16;
					out<=118;
				end
				if(in == 263) begin
					state<=16;
					out<=119;
				end
				if(in == 264) begin
					state<=16;
					out<=120;
				end
				if(in == 265) begin
					state<=16;
					out<=121;
				end
				if(in == 266) begin
					state<=16;
					out<=122;
				end
				if(in == 267) begin
					state<=16;
					out<=123;
				end
				if(in == 268) begin
					state<=16;
					out<=124;
				end
				if(in == 269) begin
					state<=16;
					out<=125;
				end
				if(in == 270) begin
					state<=16;
					out<=126;
				end
				if(in == 271) begin
					state<=16;
					out<=127;
				end
				if(in == 272) begin
					state<=16;
					out<=128;
				end
				if(in == 273) begin
					state<=16;
					out<=129;
				end
				if(in == 274) begin
					state<=16;
					out<=130;
				end
				if(in == 275) begin
					state<=16;
					out<=131;
				end
				if(in == 276) begin
					state<=16;
					out<=132;
				end
				if(in == 277) begin
					state<=16;
					out<=133;
				end
				if(in == 278) begin
					state<=16;
					out<=134;
				end
				if(in == 279) begin
					state<=16;
					out<=135;
				end
				if(in == 280) begin
					state<=16;
					out<=136;
				end
				if(in == 281) begin
					state<=16;
					out<=137;
				end
				if(in == 282) begin
					state<=16;
					out<=138;
				end
				if(in == 283) begin
					state<=16;
					out<=139;
				end
				if(in == 284) begin
					state<=16;
					out<=140;
				end
				if(in == 285) begin
					state<=16;
					out<=141;
				end
				if(in == 286) begin
					state<=16;
					out<=142;
				end
				if(in == 287) begin
					state<=16;
					out<=143;
				end
				if(in == 288) begin
					state<=16;
					out<=144;
				end
				if(in == 289) begin
					state<=16;
					out<=145;
				end
				if(in == 290) begin
					state<=16;
					out<=146;
				end
				if(in == 291) begin
					state<=16;
					out<=147;
				end
				if(in == 292) begin
					state<=16;
					out<=148;
				end
				if(in == 293) begin
					state<=16;
					out<=149;
				end
				if(in == 294) begin
					state<=16;
					out<=150;
				end
				if(in == 295) begin
					state<=16;
					out<=151;
				end
				if(in == 296) begin
					state<=16;
					out<=152;
				end
				if(in == 297) begin
					state<=16;
					out<=153;
				end
				if(in == 298) begin
					state<=16;
					out<=154;
				end
				if(in == 299) begin
					state<=16;
					out<=155;
				end
				if(in == 300) begin
					state<=16;
					out<=156;
				end
				if(in == 301) begin
					state<=16;
					out<=157;
				end
				if(in == 302) begin
					state<=16;
					out<=158;
				end
				if(in == 303) begin
					state<=16;
					out<=159;
				end
				if(in == 304) begin
					state<=16;
					out<=160;
				end
				if(in == 305) begin
					state<=16;
					out<=161;
				end
				if(in == 306) begin
					state<=16;
					out<=162;
				end
				if(in == 307) begin
					state<=16;
					out<=163;
				end
				if(in == 308) begin
					state<=16;
					out<=164;
				end
				if(in == 309) begin
					state<=16;
					out<=165;
				end
				if(in == 310) begin
					state<=16;
					out<=166;
				end
				if(in == 311) begin
					state<=16;
					out<=167;
				end
				if(in == 312) begin
					state<=16;
					out<=168;
				end
				if(in == 313) begin
					state<=16;
					out<=169;
				end
				if(in == 314) begin
					state<=16;
					out<=170;
				end
				if(in == 315) begin
					state<=16;
					out<=171;
				end
				if(in == 316) begin
					state<=16;
					out<=172;
				end
				if(in == 317) begin
					state<=16;
					out<=173;
				end
				if(in == 318) begin
					state<=16;
					out<=174;
				end
				if(in == 319) begin
					state<=16;
					out<=175;
				end
				if(in == 320) begin
					state<=16;
					out<=176;
				end
				if(in == 321) begin
					state<=16;
					out<=177;
				end
				if(in == 322) begin
					state<=16;
					out<=178;
				end
				if(in == 323) begin
					state<=16;
					out<=179;
				end
				if(in == 324) begin
					state<=16;
					out<=180;
				end
				if(in == 325) begin
					state<=16;
					out<=181;
				end
				if(in == 326) begin
					state<=16;
					out<=182;
				end
				if(in == 327) begin
					state<=16;
					out<=183;
				end
				if(in == 328) begin
					state<=16;
					out<=184;
				end
				if(in == 329) begin
					state<=16;
					out<=185;
				end
				if(in == 330) begin
					state<=16;
					out<=186;
				end
				if(in == 331) begin
					state<=16;
					out<=187;
				end
				if(in == 332) begin
					state<=16;
					out<=188;
				end
				if(in == 333) begin
					state<=16;
					out<=189;
				end
				if(in == 334) begin
					state<=16;
					out<=190;
				end
				if(in == 335) begin
					state<=16;
					out<=191;
				end
				if(in == 336) begin
					state<=16;
					out<=192;
				end
				if(in == 337) begin
					state<=16;
					out<=193;
				end
				if(in == 338) begin
					state<=16;
					out<=194;
				end
				if(in == 339) begin
					state<=16;
					out<=195;
				end
				if(in == 340) begin
					state<=16;
					out<=196;
				end
				if(in == 341) begin
					state<=16;
					out<=197;
				end
				if(in == 342) begin
					state<=16;
					out<=198;
				end
				if(in == 343) begin
					state<=16;
					out<=199;
				end
				if(in == 344) begin
					state<=16;
					out<=200;
				end
				if(in == 345) begin
					state<=16;
					out<=201;
				end
				if(in == 346) begin
					state<=16;
					out<=202;
				end
				if(in == 347) begin
					state<=16;
					out<=203;
				end
				if(in == 348) begin
					state<=16;
					out<=204;
				end
				if(in == 349) begin
					state<=16;
					out<=205;
				end
				if(in == 350) begin
					state<=16;
					out<=206;
				end
				if(in == 351) begin
					state<=16;
					out<=207;
				end
				if(in == 352) begin
					state<=16;
					out<=208;
				end
				if(in == 353) begin
					state<=16;
					out<=209;
				end
				if(in == 354) begin
					state<=16;
					out<=210;
				end
				if(in == 355) begin
					state<=16;
					out<=211;
				end
				if(in == 356) begin
					state<=16;
					out<=212;
				end
				if(in == 357) begin
					state<=16;
					out<=213;
				end
				if(in == 358) begin
					state<=16;
					out<=214;
				end
				if(in == 359) begin
					state<=16;
					out<=215;
				end
				if(in == 360) begin
					state<=16;
					out<=216;
				end
				if(in == 361) begin
					state<=16;
					out<=217;
				end
				if(in == 362) begin
					state<=16;
					out<=218;
				end
				if(in == 363) begin
					state<=16;
					out<=219;
				end
				if(in == 364) begin
					state<=16;
					out<=220;
				end
				if(in == 365) begin
					state<=16;
					out<=221;
				end
				if(in == 366) begin
					state<=16;
					out<=222;
				end
				if(in == 367) begin
					state<=16;
					out<=223;
				end
				if(in == 368) begin
					state<=16;
					out<=224;
				end
				if(in == 369) begin
					state<=16;
					out<=225;
				end
				if(in == 370) begin
					state<=16;
					out<=226;
				end
				if(in == 371) begin
					state<=16;
					out<=227;
				end
				if(in == 372) begin
					state<=16;
					out<=228;
				end
				if(in == 373) begin
					state<=16;
					out<=229;
				end
				if(in == 374) begin
					state<=16;
					out<=230;
				end
				if(in == 375) begin
					state<=16;
					out<=231;
				end
				if(in == 376) begin
					state<=16;
					out<=232;
				end
				if(in == 377) begin
					state<=16;
					out<=233;
				end
				if(in == 378) begin
					state<=16;
					out<=234;
				end
				if(in == 379) begin
					state<=16;
					out<=235;
				end
				if(in == 380) begin
					state<=16;
					out<=236;
				end
				if(in == 381) begin
					state<=16;
					out<=237;
				end
				if(in == 382) begin
					state<=16;
					out<=238;
				end
				if(in == 383) begin
					state<=16;
					out<=239;
				end
				if(in == 384) begin
					state<=16;
					out<=240;
				end
				if(in == 385) begin
					state<=16;
					out<=241;
				end
				if(in == 386) begin
					state<=16;
					out<=242;
				end
				if(in == 387) begin
					state<=16;
					out<=243;
				end
				if(in == 388) begin
					state<=16;
					out<=244;
				end
				if(in == 389) begin
					state<=16;
					out<=245;
				end
				if(in == 390) begin
					state<=16;
					out<=246;
				end
				if(in == 391) begin
					state<=16;
					out<=247;
				end
				if(in == 392) begin
					state<=16;
					out<=248;
				end
				if(in == 393) begin
					state<=16;
					out<=249;
				end
				if(in == 394) begin
					state<=16;
					out<=250;
				end
				if(in == 395) begin
					state<=16;
					out<=251;
				end
				if(in == 396) begin
					state<=16;
					out<=252;
				end
				if(in == 397) begin
					state<=16;
					out<=253;
				end
				if(in == 398) begin
					state<=16;
					out<=254;
				end
				if(in == 399) begin
					state<=16;
					out<=255;
				end
				if(in == 400) begin
					state<=16;
					out<=0;
				end
				if(in == 401) begin
					state<=16;
					out<=1;
				end
				if(in == 402) begin
					state<=16;
					out<=2;
				end
				if(in == 403) begin
					state<=16;
					out<=3;
				end
				if(in == 404) begin
					state<=16;
					out<=4;
				end
				if(in == 405) begin
					state<=16;
					out<=5;
				end
				if(in == 406) begin
					state<=16;
					out<=6;
				end
				if(in == 407) begin
					state<=16;
					out<=7;
				end
				if(in == 408) begin
					state<=16;
					out<=8;
				end
				if(in == 409) begin
					state<=16;
					out<=9;
				end
				if(in == 410) begin
					state<=16;
					out<=10;
				end
				if(in == 411) begin
					state<=16;
					out<=11;
				end
				if(in == 412) begin
					state<=16;
					out<=12;
				end
				if(in == 413) begin
					state<=16;
					out<=13;
				end
				if(in == 414) begin
					state<=16;
					out<=14;
				end
				if(in == 415) begin
					state<=16;
					out<=15;
				end
				if(in == 416) begin
					state<=16;
					out<=16;
				end
				if(in == 417) begin
					state<=16;
					out<=17;
				end
				if(in == 418) begin
					state<=16;
					out<=18;
				end
				if(in == 419) begin
					state<=16;
					out<=19;
				end
				if(in == 420) begin
					state<=16;
					out<=20;
				end
				if(in == 421) begin
					state<=16;
					out<=21;
				end
				if(in == 422) begin
					state<=16;
					out<=22;
				end
				if(in == 423) begin
					state<=16;
					out<=23;
				end
				if(in == 424) begin
					state<=16;
					out<=24;
				end
				if(in == 425) begin
					state<=16;
					out<=25;
				end
				if(in == 426) begin
					state<=16;
					out<=26;
				end
				if(in == 427) begin
					state<=16;
					out<=27;
				end
				if(in == 428) begin
					state<=16;
					out<=28;
				end
				if(in == 429) begin
					state<=16;
					out<=29;
				end
				if(in == 430) begin
					state<=16;
					out<=30;
				end
				if(in == 431) begin
					state<=16;
					out<=31;
				end
				if(in == 432) begin
					state<=16;
					out<=32;
				end
				if(in == 433) begin
					state<=16;
					out<=33;
				end
				if(in == 434) begin
					state<=16;
					out<=34;
				end
				if(in == 435) begin
					state<=16;
					out<=35;
				end
				if(in == 436) begin
					state<=16;
					out<=36;
				end
				if(in == 437) begin
					state<=16;
					out<=37;
				end
				if(in == 438) begin
					state<=16;
					out<=38;
				end
				if(in == 439) begin
					state<=16;
					out<=39;
				end
				if(in == 440) begin
					state<=16;
					out<=40;
				end
				if(in == 441) begin
					state<=16;
					out<=41;
				end
				if(in == 442) begin
					state<=16;
					out<=42;
				end
				if(in == 443) begin
					state<=16;
					out<=43;
				end
				if(in == 444) begin
					state<=16;
					out<=44;
				end
				if(in == 445) begin
					state<=16;
					out<=45;
				end
				if(in == 446) begin
					state<=16;
					out<=46;
				end
				if(in == 447) begin
					state<=16;
					out<=47;
				end
				if(in == 448) begin
					state<=16;
					out<=48;
				end
				if(in == 449) begin
					state<=16;
					out<=49;
				end
				if(in == 450) begin
					state<=16;
					out<=50;
				end
				if(in == 451) begin
					state<=16;
					out<=51;
				end
				if(in == 452) begin
					state<=16;
					out<=52;
				end
				if(in == 453) begin
					state<=16;
					out<=53;
				end
				if(in == 454) begin
					state<=16;
					out<=54;
				end
				if(in == 455) begin
					state<=16;
					out<=55;
				end
				if(in == 456) begin
					state<=16;
					out<=56;
				end
				if(in == 457) begin
					state<=16;
					out<=57;
				end
				if(in == 458) begin
					state<=16;
					out<=58;
				end
				if(in == 459) begin
					state<=16;
					out<=59;
				end
				if(in == 460) begin
					state<=16;
					out<=60;
				end
				if(in == 461) begin
					state<=16;
					out<=61;
				end
				if(in == 462) begin
					state<=16;
					out<=62;
				end
				if(in == 463) begin
					state<=16;
					out<=63;
				end
				if(in == 464) begin
					state<=16;
					out<=64;
				end
				if(in == 465) begin
					state<=1;
					out<=65;
				end
				if(in == 466) begin
					state<=1;
					out<=66;
				end
				if(in == 467) begin
					state<=1;
					out<=67;
				end
				if(in == 468) begin
					state<=1;
					out<=68;
				end
				if(in == 469) begin
					state<=1;
					out<=69;
				end
				if(in == 470) begin
					state<=1;
					out<=70;
				end
				if(in == 471) begin
					state<=1;
					out<=71;
				end
				if(in == 472) begin
					state<=1;
					out<=72;
				end
				if(in == 473) begin
					state<=1;
					out<=73;
				end
				if(in == 474) begin
					state<=1;
					out<=74;
				end
				if(in == 475) begin
					state<=1;
					out<=75;
				end
				if(in == 476) begin
					state<=1;
					out<=76;
				end
				if(in == 477) begin
					state<=1;
					out<=77;
				end
				if(in == 478) begin
					state<=1;
					out<=78;
				end
				if(in == 479) begin
					state<=1;
					out<=79;
				end
				if(in == 480) begin
					state<=1;
					out<=80;
				end
				if(in == 481) begin
					state<=1;
					out<=81;
				end
				if(in == 482) begin
					state<=1;
					out<=82;
				end
				if(in == 483) begin
					state<=1;
					out<=83;
				end
				if(in == 484) begin
					state<=1;
					out<=84;
				end
				if(in == 485) begin
					state<=1;
					out<=85;
				end
				if(in == 486) begin
					state<=1;
					out<=86;
				end
				if(in == 487) begin
					state<=1;
					out<=87;
				end
				if(in == 488) begin
					state<=1;
					out<=88;
				end
				if(in == 489) begin
					state<=1;
					out<=89;
				end
				if(in == 490) begin
					state<=1;
					out<=90;
				end
				if(in == 491) begin
					state<=1;
					out<=91;
				end
				if(in == 492) begin
					state<=1;
					out<=92;
				end
				if(in == 493) begin
					state<=1;
					out<=93;
				end
				if(in == 494) begin
					state<=1;
					out<=94;
				end
				if(in == 495) begin
					state<=1;
					out<=95;
				end
				if(in == 496) begin
					state<=1;
					out<=96;
				end
				if(in == 497) begin
					state<=1;
					out<=97;
				end
				if(in == 498) begin
					state<=1;
					out<=98;
				end
				if(in == 499) begin
					state<=1;
					out<=99;
				end
				if(in == 500) begin
					state<=1;
					out<=100;
				end
				if(in == 501) begin
					state<=1;
					out<=101;
				end
				if(in == 502) begin
					state<=1;
					out<=102;
				end
				if(in == 503) begin
					state<=1;
					out<=103;
				end
				if(in == 504) begin
					state<=1;
					out<=104;
				end
				if(in == 505) begin
					state<=1;
					out<=105;
				end
				if(in == 506) begin
					state<=1;
					out<=106;
				end
				if(in == 507) begin
					state<=1;
					out<=107;
				end
				if(in == 508) begin
					state<=1;
					out<=108;
				end
				if(in == 509) begin
					state<=1;
					out<=109;
				end
				if(in == 510) begin
					state<=1;
					out<=110;
				end
				if(in == 511) begin
					state<=1;
					out<=111;
				end
				if(in == 512) begin
					state<=1;
					out<=112;
				end
				if(in == 513) begin
					state<=1;
					out<=113;
				end
				if(in == 514) begin
					state<=1;
					out<=114;
				end
				if(in == 515) begin
					state<=1;
					out<=115;
				end
				if(in == 516) begin
					state<=1;
					out<=116;
				end
				if(in == 517) begin
					state<=1;
					out<=117;
				end
				if(in == 518) begin
					state<=1;
					out<=118;
				end
				if(in == 519) begin
					state<=1;
					out<=119;
				end
				if(in == 520) begin
					state<=1;
					out<=120;
				end
				if(in == 521) begin
					state<=1;
					out<=121;
				end
				if(in == 522) begin
					state<=1;
					out<=122;
				end
				if(in == 523) begin
					state<=1;
					out<=123;
				end
				if(in == 524) begin
					state<=1;
					out<=124;
				end
				if(in == 525) begin
					state<=1;
					out<=125;
				end
				if(in == 526) begin
					state<=1;
					out<=126;
				end
				if(in == 527) begin
					state<=1;
					out<=127;
				end
				if(in == 528) begin
					state<=1;
					out<=128;
				end
				if(in == 529) begin
					state<=1;
					out<=129;
				end
				if(in == 530) begin
					state<=1;
					out<=130;
				end
				if(in == 531) begin
					state<=1;
					out<=131;
				end
				if(in == 532) begin
					state<=1;
					out<=132;
				end
				if(in == 533) begin
					state<=1;
					out<=133;
				end
				if(in == 534) begin
					state<=1;
					out<=134;
				end
				if(in == 535) begin
					state<=1;
					out<=135;
				end
				if(in == 536) begin
					state<=1;
					out<=136;
				end
				if(in == 537) begin
					state<=1;
					out<=137;
				end
				if(in == 538) begin
					state<=1;
					out<=138;
				end
				if(in == 539) begin
					state<=1;
					out<=139;
				end
				if(in == 540) begin
					state<=1;
					out<=140;
				end
				if(in == 541) begin
					state<=1;
					out<=141;
				end
				if(in == 542) begin
					state<=1;
					out<=142;
				end
				if(in == 543) begin
					state<=1;
					out<=143;
				end
				if(in == 544) begin
					state<=1;
					out<=144;
				end
				if(in == 545) begin
					state<=1;
					out<=145;
				end
				if(in == 546) begin
					state<=1;
					out<=146;
				end
				if(in == 547) begin
					state<=1;
					out<=147;
				end
				if(in == 548) begin
					state<=1;
					out<=148;
				end
				if(in == 549) begin
					state<=1;
					out<=149;
				end
				if(in == 550) begin
					state<=1;
					out<=150;
				end
				if(in == 551) begin
					state<=1;
					out<=151;
				end
				if(in == 552) begin
					state<=1;
					out<=152;
				end
				if(in == 553) begin
					state<=1;
					out<=153;
				end
				if(in == 554) begin
					state<=1;
					out<=154;
				end
				if(in == 555) begin
					state<=1;
					out<=155;
				end
				if(in == 556) begin
					state<=1;
					out<=156;
				end
				if(in == 557) begin
					state<=1;
					out<=157;
				end
				if(in == 558) begin
					state<=1;
					out<=158;
				end
				if(in == 559) begin
					state<=1;
					out<=159;
				end
				if(in == 560) begin
					state<=1;
					out<=160;
				end
				if(in == 561) begin
					state<=1;
					out<=161;
				end
				if(in == 562) begin
					state<=1;
					out<=162;
				end
				if(in == 563) begin
					state<=1;
					out<=163;
				end
				if(in == 564) begin
					state<=1;
					out<=164;
				end
				if(in == 565) begin
					state<=1;
					out<=165;
				end
				if(in == 566) begin
					state<=1;
					out<=166;
				end
				if(in == 567) begin
					state<=1;
					out<=167;
				end
				if(in == 568) begin
					state<=1;
					out<=168;
				end
				if(in == 569) begin
					state<=1;
					out<=169;
				end
				if(in == 570) begin
					state<=1;
					out<=170;
				end
				if(in == 571) begin
					state<=1;
					out<=171;
				end
				if(in == 572) begin
					state<=1;
					out<=172;
				end
				if(in == 573) begin
					state<=1;
					out<=173;
				end
				if(in == 574) begin
					state<=1;
					out<=174;
				end
				if(in == 575) begin
					state<=1;
					out<=175;
				end
				if(in == 576) begin
					state<=1;
					out<=176;
				end
				if(in == 577) begin
					state<=1;
					out<=177;
				end
				if(in == 578) begin
					state<=1;
					out<=178;
				end
				if(in == 579) begin
					state<=1;
					out<=179;
				end
				if(in == 580) begin
					state<=1;
					out<=180;
				end
				if(in == 581) begin
					state<=1;
					out<=181;
				end
				if(in == 582) begin
					state<=1;
					out<=182;
				end
				if(in == 583) begin
					state<=1;
					out<=183;
				end
				if(in == 584) begin
					state<=1;
					out<=184;
				end
				if(in == 585) begin
					state<=1;
					out<=185;
				end
				if(in == 586) begin
					state<=1;
					out<=186;
				end
				if(in == 587) begin
					state<=1;
					out<=187;
				end
				if(in == 588) begin
					state<=1;
					out<=188;
				end
				if(in == 589) begin
					state<=1;
					out<=189;
				end
				if(in == 590) begin
					state<=1;
					out<=190;
				end
				if(in == 591) begin
					state<=1;
					out<=191;
				end
				if(in == 592) begin
					state<=1;
					out<=192;
				end
				if(in == 593) begin
					state<=1;
					out<=193;
				end
				if(in == 594) begin
					state<=1;
					out<=194;
				end
				if(in == 595) begin
					state<=1;
					out<=195;
				end
				if(in == 596) begin
					state<=1;
					out<=196;
				end
				if(in == 597) begin
					state<=1;
					out<=197;
				end
				if(in == 598) begin
					state<=1;
					out<=198;
				end
				if(in == 599) begin
					state<=1;
					out<=199;
				end
				if(in == 600) begin
					state<=1;
					out<=200;
				end
				if(in == 601) begin
					state<=1;
					out<=201;
				end
				if(in == 602) begin
					state<=1;
					out<=202;
				end
				if(in == 603) begin
					state<=1;
					out<=203;
				end
				if(in == 604) begin
					state<=1;
					out<=204;
				end
				if(in == 605) begin
					state<=1;
					out<=205;
				end
				if(in == 606) begin
					state<=1;
					out<=206;
				end
				if(in == 607) begin
					state<=1;
					out<=207;
				end
				if(in == 608) begin
					state<=1;
					out<=208;
				end
				if(in == 609) begin
					state<=1;
					out<=209;
				end
				if(in == 610) begin
					state<=1;
					out<=210;
				end
				if(in == 611) begin
					state<=1;
					out<=211;
				end
				if(in == 612) begin
					state<=1;
					out<=212;
				end
				if(in == 613) begin
					state<=1;
					out<=213;
				end
				if(in == 614) begin
					state<=1;
					out<=214;
				end
				if(in == 615) begin
					state<=1;
					out<=215;
				end
				if(in == 616) begin
					state<=1;
					out<=216;
				end
				if(in == 617) begin
					state<=1;
					out<=217;
				end
				if(in == 618) begin
					state<=1;
					out<=218;
				end
				if(in == 619) begin
					state<=1;
					out<=219;
				end
				if(in == 620) begin
					state<=1;
					out<=220;
				end
				if(in == 621) begin
					state<=1;
					out<=221;
				end
				if(in == 622) begin
					state<=1;
					out<=222;
				end
				if(in == 623) begin
					state<=1;
					out<=223;
				end
				if(in == 624) begin
					state<=1;
					out<=224;
				end
				if(in == 625) begin
					state<=1;
					out<=225;
				end
				if(in == 626) begin
					state<=1;
					out<=226;
				end
				if(in == 627) begin
					state<=1;
					out<=227;
				end
				if(in == 628) begin
					state<=1;
					out<=228;
				end
				if(in == 629) begin
					state<=1;
					out<=229;
				end
				if(in == 630) begin
					state<=1;
					out<=230;
				end
				if(in == 631) begin
					state<=1;
					out<=231;
				end
				if(in == 632) begin
					state<=1;
					out<=232;
				end
				if(in == 633) begin
					state<=1;
					out<=233;
				end
				if(in == 634) begin
					state<=1;
					out<=234;
				end
				if(in == 635) begin
					state<=1;
					out<=235;
				end
				if(in == 636) begin
					state<=1;
					out<=236;
				end
				if(in == 637) begin
					state<=1;
					out<=237;
				end
				if(in == 638) begin
					state<=1;
					out<=238;
				end
				if(in == 639) begin
					state<=1;
					out<=239;
				end
				if(in == 640) begin
					state<=1;
					out<=240;
				end
				if(in == 641) begin
					state<=1;
					out<=241;
				end
				if(in == 642) begin
					state<=1;
					out<=242;
				end
				if(in == 643) begin
					state<=1;
					out<=243;
				end
				if(in == 644) begin
					state<=1;
					out<=244;
				end
				if(in == 645) begin
					state<=1;
					out<=245;
				end
				if(in == 646) begin
					state<=1;
					out<=246;
				end
				if(in == 647) begin
					state<=1;
					out<=247;
				end
				if(in == 648) begin
					state<=1;
					out<=248;
				end
				if(in == 649) begin
					state<=1;
					out<=249;
				end
				if(in == 650) begin
					state<=1;
					out<=250;
				end
				if(in == 651) begin
					state<=1;
					out<=251;
				end
				if(in == 652) begin
					state<=1;
					out<=252;
				end
				if(in == 653) begin
					state<=1;
					out<=253;
				end
				if(in == 654) begin
					state<=1;
					out<=254;
				end
				if(in == 655) begin
					state<=1;
					out<=255;
				end
				if(in == 656) begin
					state<=1;
					out<=0;
				end
				if(in == 657) begin
					state<=1;
					out<=1;
				end
				if(in == 658) begin
					state<=1;
					out<=2;
				end
				if(in == 659) begin
					state<=1;
					out<=3;
				end
				if(in == 660) begin
					state<=1;
					out<=4;
				end
				if(in == 661) begin
					state<=1;
					out<=5;
				end
				if(in == 662) begin
					state<=1;
					out<=6;
				end
				if(in == 663) begin
					state<=1;
					out<=7;
				end
				if(in == 664) begin
					state<=1;
					out<=8;
				end
				if(in == 665) begin
					state<=1;
					out<=9;
				end
				if(in == 666) begin
					state<=1;
					out<=10;
				end
				if(in == 667) begin
					state<=1;
					out<=11;
				end
				if(in == 668) begin
					state<=1;
					out<=12;
				end
				if(in == 669) begin
					state<=1;
					out<=13;
				end
				if(in == 670) begin
					state<=1;
					out<=14;
				end
				if(in == 671) begin
					state<=1;
					out<=15;
				end
				if(in == 672) begin
					state<=1;
					out<=16;
				end
				if(in == 673) begin
					state<=1;
					out<=17;
				end
				if(in == 674) begin
					state<=1;
					out<=18;
				end
				if(in == 675) begin
					state<=1;
					out<=19;
				end
				if(in == 676) begin
					state<=1;
					out<=20;
				end
				if(in == 677) begin
					state<=1;
					out<=21;
				end
				if(in == 678) begin
					state<=1;
					out<=22;
				end
				if(in == 679) begin
					state<=1;
					out<=23;
				end
				if(in == 680) begin
					state<=1;
					out<=24;
				end
				if(in == 681) begin
					state<=1;
					out<=25;
				end
				if(in == 682) begin
					state<=1;
					out<=26;
				end
				if(in == 683) begin
					state<=1;
					out<=27;
				end
				if(in == 684) begin
					state<=1;
					out<=28;
				end
				if(in == 685) begin
					state<=1;
					out<=29;
				end
				if(in == 686) begin
					state<=1;
					out<=30;
				end
				if(in == 687) begin
					state<=1;
					out<=31;
				end
				if(in == 688) begin
					state<=1;
					out<=32;
				end
				if(in == 689) begin
					state<=1;
					out<=33;
				end
				if(in == 690) begin
					state<=1;
					out<=34;
				end
				if(in == 691) begin
					state<=1;
					out<=35;
				end
				if(in == 692) begin
					state<=1;
					out<=36;
				end
				if(in == 693) begin
					state<=1;
					out<=37;
				end
				if(in == 694) begin
					state<=1;
					out<=38;
				end
				if(in == 695) begin
					state<=1;
					out<=39;
				end
				if(in == 696) begin
					state<=1;
					out<=40;
				end
				if(in == 697) begin
					state<=1;
					out<=41;
				end
				if(in == 698) begin
					state<=1;
					out<=42;
				end
				if(in == 699) begin
					state<=1;
					out<=43;
				end
				if(in == 700) begin
					state<=1;
					out<=44;
				end
				if(in == 701) begin
					state<=1;
					out<=45;
				end
				if(in == 702) begin
					state<=1;
					out<=46;
				end
				if(in == 703) begin
					state<=1;
					out<=47;
				end
				if(in == 704) begin
					state<=1;
					out<=48;
				end
				if(in == 705) begin
					state<=1;
					out<=49;
				end
				if(in == 706) begin
					state<=1;
					out<=50;
				end
				if(in == 707) begin
					state<=1;
					out<=51;
				end
				if(in == 708) begin
					state<=1;
					out<=52;
				end
				if(in == 709) begin
					state<=1;
					out<=53;
				end
				if(in == 710) begin
					state<=1;
					out<=54;
				end
				if(in == 711) begin
					state<=1;
					out<=55;
				end
				if(in == 712) begin
					state<=1;
					out<=56;
				end
				if(in == 713) begin
					state<=1;
					out<=57;
				end
				if(in == 714) begin
					state<=1;
					out<=58;
				end
				if(in == 715) begin
					state<=1;
					out<=59;
				end
				if(in == 716) begin
					state<=1;
					out<=60;
				end
				if(in == 717) begin
					state<=1;
					out<=61;
				end
				if(in == 718) begin
					state<=1;
					out<=62;
				end
				if(in == 719) begin
					state<=1;
					out<=63;
				end
				if(in == 720) begin
					state<=1;
					out<=64;
				end
				if(in == 721) begin
					state<=1;
					out<=65;
				end
				if(in == 722) begin
					state<=1;
					out<=66;
				end
				if(in == 723) begin
					state<=1;
					out<=67;
				end
				if(in == 724) begin
					state<=1;
					out<=68;
				end
				if(in == 725) begin
					state<=1;
					out<=69;
				end
				if(in == 726) begin
					state<=1;
					out<=70;
				end
				if(in == 727) begin
					state<=1;
					out<=71;
				end
				if(in == 728) begin
					state<=1;
					out<=72;
				end
				if(in == 729) begin
					state<=1;
					out<=73;
				end
				if(in == 730) begin
					state<=1;
					out<=74;
				end
				if(in == 731) begin
					state<=1;
					out<=75;
				end
				if(in == 732) begin
					state<=1;
					out<=76;
				end
				if(in == 733) begin
					state<=1;
					out<=77;
				end
				if(in == 734) begin
					state<=1;
					out<=78;
				end
				if(in == 735) begin
					state<=1;
					out<=79;
				end
				if(in == 736) begin
					state<=1;
					out<=80;
				end
				if(in == 737) begin
					state<=1;
					out<=81;
				end
				if(in == 738) begin
					state<=1;
					out<=82;
				end
				if(in == 739) begin
					state<=1;
					out<=83;
				end
				if(in == 740) begin
					state<=1;
					out<=84;
				end
				if(in == 741) begin
					state<=1;
					out<=85;
				end
				if(in == 742) begin
					state<=1;
					out<=86;
				end
				if(in == 743) begin
					state<=1;
					out<=87;
				end
				if(in == 744) begin
					state<=1;
					out<=88;
				end
				if(in == 745) begin
					state<=1;
					out<=89;
				end
				if(in == 746) begin
					state<=1;
					out<=90;
				end
				if(in == 747) begin
					state<=1;
					out<=91;
				end
				if(in == 748) begin
					state<=1;
					out<=92;
				end
				if(in == 749) begin
					state<=1;
					out<=93;
				end
				if(in == 750) begin
					state<=1;
					out<=94;
				end
				if(in == 751) begin
					state<=1;
					out<=95;
				end
				if(in == 752) begin
					state<=1;
					out<=96;
				end
				if(in == 753) begin
					state<=1;
					out<=97;
				end
				if(in == 754) begin
					state<=1;
					out<=98;
				end
				if(in == 755) begin
					state<=1;
					out<=99;
				end
				if(in == 756) begin
					state<=1;
					out<=100;
				end
				if(in == 757) begin
					state<=1;
					out<=101;
				end
				if(in == 758) begin
					state<=1;
					out<=102;
				end
				if(in == 759) begin
					state<=1;
					out<=103;
				end
				if(in == 760) begin
					state<=1;
					out<=104;
				end
				if(in == 761) begin
					state<=1;
					out<=105;
				end
				if(in == 762) begin
					state<=1;
					out<=106;
				end
				if(in == 763) begin
					state<=1;
					out<=107;
				end
				if(in == 764) begin
					state<=1;
					out<=108;
				end
				if(in == 765) begin
					state<=1;
					out<=109;
				end
				if(in == 766) begin
					state<=1;
					out<=110;
				end
				if(in == 767) begin
					state<=1;
					out<=111;
				end
				if(in == 768) begin
					state<=1;
					out<=112;
				end
				if(in == 769) begin
					state<=1;
					out<=113;
				end
				if(in == 770) begin
					state<=1;
					out<=114;
				end
				if(in == 771) begin
					state<=1;
					out<=115;
				end
				if(in == 772) begin
					state<=1;
					out<=116;
				end
				if(in == 773) begin
					state<=1;
					out<=117;
				end
				if(in == 774) begin
					state<=1;
					out<=118;
				end
				if(in == 775) begin
					state<=1;
					out<=119;
				end
				if(in == 776) begin
					state<=1;
					out<=120;
				end
				if(in == 777) begin
					state<=1;
					out<=121;
				end
				if(in == 778) begin
					state<=1;
					out<=122;
				end
				if(in == 779) begin
					state<=1;
					out<=123;
				end
				if(in == 780) begin
					state<=1;
					out<=124;
				end
				if(in == 781) begin
					state<=1;
					out<=125;
				end
				if(in == 782) begin
					state<=1;
					out<=126;
				end
				if(in == 783) begin
					state<=1;
					out<=127;
				end
				if(in == 784) begin
					state<=1;
					out<=128;
				end
				if(in == 785) begin
					state<=1;
					out<=129;
				end
				if(in == 786) begin
					state<=1;
					out<=130;
				end
				if(in == 787) begin
					state<=1;
					out<=131;
				end
				if(in == 788) begin
					state<=1;
					out<=132;
				end
				if(in == 789) begin
					state<=1;
					out<=133;
				end
				if(in == 790) begin
					state<=1;
					out<=134;
				end
				if(in == 791) begin
					state<=1;
					out<=135;
				end
				if(in == 792) begin
					state<=1;
					out<=136;
				end
				if(in == 793) begin
					state<=1;
					out<=137;
				end
				if(in == 794) begin
					state<=1;
					out<=138;
				end
				if(in == 795) begin
					state<=1;
					out<=139;
				end
				if(in == 796) begin
					state<=1;
					out<=140;
				end
				if(in == 797) begin
					state<=1;
					out<=141;
				end
				if(in == 798) begin
					state<=1;
					out<=142;
				end
				if(in == 799) begin
					state<=1;
					out<=143;
				end
				if(in == 800) begin
					state<=1;
					out<=144;
				end
				if(in == 801) begin
					state<=1;
					out<=145;
				end
				if(in == 802) begin
					state<=1;
					out<=146;
				end
				if(in == 803) begin
					state<=1;
					out<=147;
				end
				if(in == 804) begin
					state<=1;
					out<=148;
				end
				if(in == 805) begin
					state<=1;
					out<=149;
				end
				if(in == 806) begin
					state<=1;
					out<=150;
				end
				if(in == 807) begin
					state<=1;
					out<=151;
				end
				if(in == 808) begin
					state<=1;
					out<=152;
				end
				if(in == 809) begin
					state<=1;
					out<=153;
				end
				if(in == 810) begin
					state<=1;
					out<=154;
				end
				if(in == 811) begin
					state<=1;
					out<=155;
				end
				if(in == 812) begin
					state<=1;
					out<=156;
				end
				if(in == 813) begin
					state<=1;
					out<=157;
				end
				if(in == 814) begin
					state<=1;
					out<=158;
				end
				if(in == 815) begin
					state<=1;
					out<=159;
				end
				if(in == 816) begin
					state<=1;
					out<=160;
				end
				if(in == 817) begin
					state<=1;
					out<=161;
				end
				if(in == 818) begin
					state<=1;
					out<=162;
				end
				if(in == 819) begin
					state<=1;
					out<=163;
				end
				if(in == 820) begin
					state<=1;
					out<=164;
				end
				if(in == 821) begin
					state<=1;
					out<=165;
				end
				if(in == 822) begin
					state<=1;
					out<=166;
				end
				if(in == 823) begin
					state<=1;
					out<=167;
				end
				if(in == 824) begin
					state<=1;
					out<=168;
				end
				if(in == 825) begin
					state<=1;
					out<=169;
				end
				if(in == 826) begin
					state<=1;
					out<=170;
				end
				if(in == 827) begin
					state<=1;
					out<=171;
				end
				if(in == 828) begin
					state<=1;
					out<=172;
				end
				if(in == 829) begin
					state<=1;
					out<=173;
				end
				if(in == 830) begin
					state<=1;
					out<=174;
				end
				if(in == 831) begin
					state<=1;
					out<=175;
				end
				if(in == 832) begin
					state<=1;
					out<=176;
				end
				if(in == 833) begin
					state<=1;
					out<=177;
				end
				if(in == 834) begin
					state<=1;
					out<=178;
				end
				if(in == 835) begin
					state<=1;
					out<=179;
				end
				if(in == 836) begin
					state<=1;
					out<=180;
				end
				if(in == 837) begin
					state<=1;
					out<=181;
				end
				if(in == 838) begin
					state<=1;
					out<=182;
				end
				if(in == 839) begin
					state<=1;
					out<=183;
				end
				if(in == 840) begin
					state<=1;
					out<=184;
				end
				if(in == 841) begin
					state<=1;
					out<=185;
				end
				if(in == 842) begin
					state<=1;
					out<=186;
				end
				if(in == 843) begin
					state<=1;
					out<=187;
				end
				if(in == 844) begin
					state<=1;
					out<=188;
				end
				if(in == 845) begin
					state<=1;
					out<=189;
				end
				if(in == 846) begin
					state<=1;
					out<=190;
				end
				if(in == 847) begin
					state<=1;
					out<=191;
				end
				if(in == 848) begin
					state<=1;
					out<=192;
				end
				if(in == 849) begin
					state<=1;
					out<=193;
				end
				if(in == 850) begin
					state<=1;
					out<=194;
				end
				if(in == 851) begin
					state<=1;
					out<=195;
				end
				if(in == 852) begin
					state<=1;
					out<=196;
				end
				if(in == 853) begin
					state<=1;
					out<=197;
				end
				if(in == 854) begin
					state<=1;
					out<=198;
				end
				if(in == 855) begin
					state<=1;
					out<=199;
				end
				if(in == 856) begin
					state<=1;
					out<=200;
				end
				if(in == 857) begin
					state<=1;
					out<=201;
				end
				if(in == 858) begin
					state<=1;
					out<=202;
				end
				if(in == 859) begin
					state<=1;
					out<=203;
				end
				if(in == 860) begin
					state<=1;
					out<=204;
				end
				if(in == 861) begin
					state<=1;
					out<=205;
				end
				if(in == 862) begin
					state<=1;
					out<=206;
				end
				if(in == 863) begin
					state<=1;
					out<=207;
				end
				if(in == 864) begin
					state<=1;
					out<=208;
				end
				if(in == 865) begin
					state<=1;
					out<=209;
				end
				if(in == 866) begin
					state<=1;
					out<=210;
				end
				if(in == 867) begin
					state<=1;
					out<=211;
				end
				if(in == 868) begin
					state<=1;
					out<=212;
				end
				if(in == 869) begin
					state<=1;
					out<=213;
				end
				if(in == 870) begin
					state<=1;
					out<=214;
				end
				if(in == 871) begin
					state<=1;
					out<=215;
				end
				if(in == 872) begin
					state<=1;
					out<=216;
				end
				if(in == 873) begin
					state<=1;
					out<=217;
				end
				if(in == 874) begin
					state<=1;
					out<=218;
				end
				if(in == 875) begin
					state<=1;
					out<=219;
				end
				if(in == 876) begin
					state<=1;
					out<=220;
				end
				if(in == 877) begin
					state<=1;
					out<=221;
				end
				if(in == 878) begin
					state<=1;
					out<=222;
				end
				if(in == 879) begin
					state<=1;
					out<=223;
				end
				if(in == 880) begin
					state<=1;
					out<=224;
				end
				if(in == 881) begin
					state<=1;
					out<=225;
				end
				if(in == 882) begin
					state<=1;
					out<=226;
				end
				if(in == 883) begin
					state<=1;
					out<=227;
				end
				if(in == 884) begin
					state<=1;
					out<=228;
				end
				if(in == 885) begin
					state<=1;
					out<=229;
				end
				if(in == 886) begin
					state<=1;
					out<=230;
				end
				if(in == 887) begin
					state<=1;
					out<=231;
				end
				if(in == 888) begin
					state<=1;
					out<=232;
				end
				if(in == 889) begin
					state<=1;
					out<=233;
				end
				if(in == 890) begin
					state<=1;
					out<=234;
				end
				if(in == 891) begin
					state<=1;
					out<=235;
				end
				if(in == 892) begin
					state<=1;
					out<=236;
				end
				if(in == 893) begin
					state<=1;
					out<=237;
				end
				if(in == 894) begin
					state<=1;
					out<=238;
				end
				if(in == 895) begin
					state<=1;
					out<=239;
				end
				if(in == 896) begin
					state<=1;
					out<=240;
				end
				if(in == 897) begin
					state<=1;
					out<=241;
				end
				if(in == 898) begin
					state<=1;
					out<=242;
				end
				if(in == 899) begin
					state<=1;
					out<=243;
				end
				if(in == 900) begin
					state<=1;
					out<=244;
				end
				if(in == 901) begin
					state<=1;
					out<=245;
				end
				if(in == 902) begin
					state<=1;
					out<=246;
				end
				if(in == 903) begin
					state<=1;
					out<=247;
				end
				if(in == 904) begin
					state<=1;
					out<=248;
				end
				if(in == 905) begin
					state<=1;
					out<=249;
				end
				if(in == 906) begin
					state<=1;
					out<=250;
				end
				if(in == 907) begin
					state<=1;
					out<=251;
				end
				if(in == 908) begin
					state<=1;
					out<=252;
				end
				if(in == 909) begin
					state<=1;
					out<=253;
				end
				if(in == 910) begin
					state<=1;
					out<=254;
				end
				if(in == 911) begin
					state<=1;
					out<=255;
				end
				if(in == 912) begin
					state<=1;
					out<=0;
				end
				if(in == 913) begin
					state<=1;
					out<=1;
				end
				if(in == 914) begin
					state<=1;
					out<=2;
				end
				if(in == 915) begin
					state<=1;
					out<=3;
				end
				if(in == 916) begin
					state<=1;
					out<=4;
				end
				if(in == 917) begin
					state<=1;
					out<=5;
				end
				if(in == 918) begin
					state<=1;
					out<=6;
				end
				if(in == 919) begin
					state<=1;
					out<=7;
				end
				if(in == 920) begin
					state<=1;
					out<=8;
				end
				if(in == 921) begin
					state<=1;
					out<=9;
				end
				if(in == 922) begin
					state<=1;
					out<=10;
				end
				if(in == 923) begin
					state<=1;
					out<=11;
				end
				if(in == 924) begin
					state<=1;
					out<=12;
				end
				if(in == 925) begin
					state<=1;
					out<=13;
				end
				if(in == 926) begin
					state<=1;
					out<=14;
				end
				if(in == 927) begin
					state<=1;
					out<=15;
				end
				if(in == 928) begin
					state<=1;
					out<=16;
				end
			end
			17: begin
				if(in == 0) begin
					state<=1;
					out<=17;
				end
				if(in == 1) begin
					state<=1;
					out<=18;
				end
				if(in == 2) begin
					state<=17;
					out<=19;
				end
				if(in == 3) begin
					state<=1;
					out<=20;
				end
				if(in == 4) begin
					state<=17;
					out<=21;
				end
				if(in == 5) begin
					state<=1;
					out<=22;
				end
				if(in == 6) begin
					state<=17;
					out<=23;
				end
				if(in == 7) begin
					state<=17;
					out<=24;
				end
				if(in == 8) begin
					state<=17;
					out<=25;
				end
				if(in == 9) begin
					state<=17;
					out<=26;
				end
				if(in == 10) begin
					state<=17;
					out<=27;
				end
				if(in == 11) begin
					state<=17;
					out<=28;
				end
				if(in == 12) begin
					state<=17;
					out<=29;
				end
				if(in == 13) begin
					state<=17;
					out<=30;
				end
				if(in == 14) begin
					state<=17;
					out<=31;
				end
				if(in == 15) begin
					state<=17;
					out<=32;
				end
				if(in == 16) begin
					state<=17;
					out<=33;
				end
				if(in == 17) begin
					state<=17;
					out<=34;
				end
				if(in == 18) begin
					state<=17;
					out<=35;
				end
				if(in == 19) begin
					state<=17;
					out<=36;
				end
				if(in == 20) begin
					state<=17;
					out<=37;
				end
				if(in == 21) begin
					state<=17;
					out<=38;
				end
				if(in == 22) begin
					state<=17;
					out<=39;
				end
				if(in == 23) begin
					state<=17;
					out<=40;
				end
				if(in == 24) begin
					state<=17;
					out<=41;
				end
				if(in == 25) begin
					state<=17;
					out<=42;
				end
				if(in == 26) begin
					state<=17;
					out<=43;
				end
				if(in == 27) begin
					state<=17;
					out<=44;
				end
				if(in == 28) begin
					state<=17;
					out<=45;
				end
				if(in == 29) begin
					state<=17;
					out<=46;
				end
				if(in == 30) begin
					state<=17;
					out<=47;
				end
				if(in == 31) begin
					state<=17;
					out<=48;
				end
				if(in == 32) begin
					state<=17;
					out<=49;
				end
				if(in == 33) begin
					state<=17;
					out<=50;
				end
				if(in == 34) begin
					state<=17;
					out<=51;
				end
				if(in == 35) begin
					state<=17;
					out<=52;
				end
				if(in == 36) begin
					state<=17;
					out<=53;
				end
				if(in == 37) begin
					state<=17;
					out<=54;
				end
				if(in == 38) begin
					state<=17;
					out<=55;
				end
				if(in == 39) begin
					state<=17;
					out<=56;
				end
				if(in == 40) begin
					state<=17;
					out<=57;
				end
				if(in == 41) begin
					state<=17;
					out<=58;
				end
				if(in == 42) begin
					state<=17;
					out<=59;
				end
				if(in == 43) begin
					state<=17;
					out<=60;
				end
				if(in == 44) begin
					state<=17;
					out<=61;
				end
				if(in == 45) begin
					state<=17;
					out<=62;
				end
				if(in == 46) begin
					state<=17;
					out<=63;
				end
				if(in == 47) begin
					state<=17;
					out<=64;
				end
				if(in == 48) begin
					state<=17;
					out<=65;
				end
				if(in == 49) begin
					state<=17;
					out<=66;
				end
				if(in == 50) begin
					state<=17;
					out<=67;
				end
				if(in == 51) begin
					state<=17;
					out<=68;
				end
				if(in == 52) begin
					state<=17;
					out<=69;
				end
				if(in == 53) begin
					state<=1;
					out<=70;
				end
				if(in == 54) begin
					state<=17;
					out<=71;
				end
				if(in == 55) begin
					state<=1;
					out<=72;
				end
				if(in == 56) begin
					state<=17;
					out<=73;
				end
				if(in == 57) begin
					state<=1;
					out<=74;
				end
				if(in == 58) begin
					state<=17;
					out<=75;
				end
				if(in == 59) begin
					state<=17;
					out<=76;
				end
				if(in == 60) begin
					state<=17;
					out<=77;
				end
				if(in == 61) begin
					state<=17;
					out<=78;
				end
				if(in == 62) begin
					state<=17;
					out<=79;
				end
				if(in == 63) begin
					state<=17;
					out<=80;
				end
				if(in == 64) begin
					state<=17;
					out<=81;
				end
				if(in == 65) begin
					state<=17;
					out<=82;
				end
				if(in == 66) begin
					state<=17;
					out<=83;
				end
				if(in == 67) begin
					state<=17;
					out<=84;
				end
				if(in == 68) begin
					state<=17;
					out<=85;
				end
				if(in == 69) begin
					state<=17;
					out<=86;
				end
				if(in == 70) begin
					state<=17;
					out<=87;
				end
				if(in == 71) begin
					state<=17;
					out<=88;
				end
				if(in == 72) begin
					state<=17;
					out<=89;
				end
				if(in == 73) begin
					state<=17;
					out<=90;
				end
				if(in == 74) begin
					state<=17;
					out<=91;
				end
				if(in == 75) begin
					state<=17;
					out<=92;
				end
				if(in == 76) begin
					state<=17;
					out<=93;
				end
				if(in == 77) begin
					state<=17;
					out<=94;
				end
				if(in == 78) begin
					state<=17;
					out<=95;
				end
				if(in == 79) begin
					state<=17;
					out<=96;
				end
				if(in == 80) begin
					state<=17;
					out<=97;
				end
				if(in == 81) begin
					state<=17;
					out<=98;
				end
				if(in == 82) begin
					state<=17;
					out<=99;
				end
				if(in == 83) begin
					state<=17;
					out<=100;
				end
				if(in == 84) begin
					state<=17;
					out<=101;
				end
				if(in == 85) begin
					state<=17;
					out<=102;
				end
				if(in == 86) begin
					state<=17;
					out<=103;
				end
				if(in == 87) begin
					state<=17;
					out<=104;
				end
				if(in == 88) begin
					state<=17;
					out<=105;
				end
				if(in == 89) begin
					state<=17;
					out<=106;
				end
				if(in == 90) begin
					state<=17;
					out<=107;
				end
				if(in == 91) begin
					state<=17;
					out<=108;
				end
				if(in == 92) begin
					state<=17;
					out<=109;
				end
				if(in == 93) begin
					state<=17;
					out<=110;
				end
				if(in == 94) begin
					state<=17;
					out<=111;
				end
				if(in == 95) begin
					state<=17;
					out<=112;
				end
				if(in == 96) begin
					state<=17;
					out<=113;
				end
				if(in == 97) begin
					state<=17;
					out<=114;
				end
				if(in == 98) begin
					state<=17;
					out<=115;
				end
				if(in == 99) begin
					state<=17;
					out<=116;
				end
				if(in == 100) begin
					state<=17;
					out<=117;
				end
				if(in == 101) begin
					state<=17;
					out<=118;
				end
				if(in == 102) begin
					state<=17;
					out<=119;
				end
				if(in == 103) begin
					state<=17;
					out<=120;
				end
				if(in == 104) begin
					state<=17;
					out<=121;
				end
				if(in == 105) begin
					state<=1;
					out<=122;
				end
				if(in == 106) begin
					state<=17;
					out<=123;
				end
				if(in == 107) begin
					state<=1;
					out<=124;
				end
				if(in == 108) begin
					state<=17;
					out<=125;
				end
				if(in == 109) begin
					state<=1;
					out<=126;
				end
				if(in == 110) begin
					state<=17;
					out<=127;
				end
				if(in == 111) begin
					state<=1;
					out<=128;
				end
				if(in == 112) begin
					state<=17;
					out<=129;
				end
				if(in == 113) begin
					state<=1;
					out<=130;
				end
				if(in == 114) begin
					state<=17;
					out<=131;
				end
				if(in == 115) begin
					state<=1;
					out<=132;
				end
				if(in == 116) begin
					state<=17;
					out<=133;
				end
				if(in == 117) begin
					state<=1;
					out<=134;
				end
				if(in == 118) begin
					state<=17;
					out<=135;
				end
				if(in == 119) begin
					state<=1;
					out<=136;
				end
				if(in == 120) begin
					state<=17;
					out<=137;
				end
				if(in == 121) begin
					state<=1;
					out<=138;
				end
				if(in == 122) begin
					state<=17;
					out<=139;
				end
				if(in == 123) begin
					state<=17;
					out<=140;
				end
				if(in == 124) begin
					state<=17;
					out<=141;
				end
				if(in == 125) begin
					state<=17;
					out<=142;
				end
				if(in == 126) begin
					state<=17;
					out<=143;
				end
				if(in == 127) begin
					state<=17;
					out<=144;
				end
				if(in == 128) begin
					state<=17;
					out<=145;
				end
				if(in == 129) begin
					state<=17;
					out<=146;
				end
				if(in == 130) begin
					state<=17;
					out<=147;
				end
				if(in == 131) begin
					state<=17;
					out<=148;
				end
				if(in == 132) begin
					state<=17;
					out<=149;
				end
				if(in == 133) begin
					state<=17;
					out<=150;
				end
				if(in == 134) begin
					state<=17;
					out<=151;
				end
				if(in == 135) begin
					state<=17;
					out<=152;
				end
				if(in == 136) begin
					state<=17;
					out<=153;
				end
				if(in == 137) begin
					state<=17;
					out<=154;
				end
				if(in == 138) begin
					state<=17;
					out<=155;
				end
				if(in == 139) begin
					state<=17;
					out<=156;
				end
				if(in == 140) begin
					state<=17;
					out<=157;
				end
				if(in == 141) begin
					state<=17;
					out<=158;
				end
				if(in == 142) begin
					state<=17;
					out<=159;
				end
				if(in == 143) begin
					state<=17;
					out<=160;
				end
				if(in == 144) begin
					state<=17;
					out<=161;
				end
				if(in == 145) begin
					state<=17;
					out<=162;
				end
				if(in == 146) begin
					state<=17;
					out<=163;
				end
				if(in == 147) begin
					state<=17;
					out<=164;
				end
				if(in == 148) begin
					state<=17;
					out<=165;
				end
				if(in == 149) begin
					state<=17;
					out<=166;
				end
				if(in == 150) begin
					state<=17;
					out<=167;
				end
				if(in == 151) begin
					state<=17;
					out<=168;
				end
				if(in == 152) begin
					state<=17;
					out<=169;
				end
				if(in == 153) begin
					state<=17;
					out<=170;
				end
				if(in == 154) begin
					state<=17;
					out<=171;
				end
				if(in == 155) begin
					state<=17;
					out<=172;
				end
				if(in == 156) begin
					state<=17;
					out<=173;
				end
				if(in == 157) begin
					state<=17;
					out<=174;
				end
				if(in == 158) begin
					state<=17;
					out<=175;
				end
				if(in == 159) begin
					state<=17;
					out<=176;
				end
				if(in == 160) begin
					state<=17;
					out<=177;
				end
				if(in == 161) begin
					state<=17;
					out<=178;
				end
				if(in == 162) begin
					state<=17;
					out<=179;
				end
				if(in == 163) begin
					state<=17;
					out<=180;
				end
				if(in == 164) begin
					state<=17;
					out<=181;
				end
				if(in == 165) begin
					state<=17;
					out<=182;
				end
				if(in == 166) begin
					state<=17;
					out<=183;
				end
				if(in == 167) begin
					state<=17;
					out<=184;
				end
				if(in == 168) begin
					state<=17;
					out<=185;
				end
				if(in == 169) begin
					state<=1;
					out<=186;
				end
				if(in == 170) begin
					state<=17;
					out<=187;
				end
				if(in == 171) begin
					state<=1;
					out<=188;
				end
				if(in == 172) begin
					state<=17;
					out<=189;
				end
				if(in == 173) begin
					state<=1;
					out<=190;
				end
				if(in == 174) begin
					state<=17;
					out<=191;
				end
				if(in == 175) begin
					state<=17;
					out<=192;
				end
				if(in == 176) begin
					state<=17;
					out<=193;
				end
				if(in == 177) begin
					state<=17;
					out<=194;
				end
				if(in == 178) begin
					state<=17;
					out<=195;
				end
				if(in == 179) begin
					state<=17;
					out<=196;
				end
				if(in == 180) begin
					state<=17;
					out<=197;
				end
				if(in == 181) begin
					state<=17;
					out<=198;
				end
				if(in == 182) begin
					state<=17;
					out<=199;
				end
				if(in == 183) begin
					state<=17;
					out<=200;
				end
				if(in == 184) begin
					state<=17;
					out<=201;
				end
				if(in == 185) begin
					state<=17;
					out<=202;
				end
				if(in == 186) begin
					state<=17;
					out<=203;
				end
				if(in == 187) begin
					state<=17;
					out<=204;
				end
				if(in == 188) begin
					state<=17;
					out<=205;
				end
				if(in == 189) begin
					state<=17;
					out<=206;
				end
				if(in == 190) begin
					state<=17;
					out<=207;
				end
				if(in == 191) begin
					state<=17;
					out<=208;
				end
				if(in == 192) begin
					state<=17;
					out<=209;
				end
				if(in == 193) begin
					state<=17;
					out<=210;
				end
				if(in == 194) begin
					state<=17;
					out<=211;
				end
				if(in == 195) begin
					state<=17;
					out<=212;
				end
				if(in == 196) begin
					state<=17;
					out<=213;
				end
				if(in == 197) begin
					state<=17;
					out<=214;
				end
				if(in == 198) begin
					state<=17;
					out<=215;
				end
				if(in == 199) begin
					state<=17;
					out<=216;
				end
				if(in == 200) begin
					state<=17;
					out<=217;
				end
				if(in == 201) begin
					state<=17;
					out<=218;
				end
				if(in == 202) begin
					state<=17;
					out<=219;
				end
				if(in == 203) begin
					state<=17;
					out<=220;
				end
				if(in == 204) begin
					state<=17;
					out<=221;
				end
				if(in == 205) begin
					state<=17;
					out<=222;
				end
				if(in == 206) begin
					state<=17;
					out<=223;
				end
				if(in == 207) begin
					state<=17;
					out<=224;
				end
				if(in == 208) begin
					state<=17;
					out<=225;
				end
				if(in == 209) begin
					state<=17;
					out<=226;
				end
				if(in == 210) begin
					state<=17;
					out<=227;
				end
				if(in == 211) begin
					state<=17;
					out<=228;
				end
				if(in == 212) begin
					state<=17;
					out<=229;
				end
				if(in == 213) begin
					state<=17;
					out<=230;
				end
				if(in == 214) begin
					state<=17;
					out<=231;
				end
				if(in == 215) begin
					state<=17;
					out<=232;
				end
				if(in == 216) begin
					state<=17;
					out<=233;
				end
				if(in == 217) begin
					state<=17;
					out<=234;
				end
				if(in == 218) begin
					state<=17;
					out<=235;
				end
				if(in == 219) begin
					state<=17;
					out<=236;
				end
				if(in == 220) begin
					state<=17;
					out<=237;
				end
				if(in == 221) begin
					state<=1;
					out<=238;
				end
				if(in == 222) begin
					state<=17;
					out<=239;
				end
				if(in == 223) begin
					state<=1;
					out<=240;
				end
				if(in == 224) begin
					state<=17;
					out<=241;
				end
				if(in == 225) begin
					state<=1;
					out<=242;
				end
				if(in == 226) begin
					state<=17;
					out<=243;
				end
				if(in == 227) begin
					state<=1;
					out<=244;
				end
				if(in == 228) begin
					state<=17;
					out<=245;
				end
				if(in == 229) begin
					state<=1;
					out<=246;
				end
				if(in == 230) begin
					state<=17;
					out<=247;
				end
				if(in == 231) begin
					state<=1;
					out<=248;
				end
				if(in == 232) begin
					state<=17;
					out<=249;
				end
				if(in == 233) begin
					state<=1;
					out<=250;
				end
				if(in == 234) begin
					state<=17;
					out<=251;
				end
				if(in == 235) begin
					state<=1;
					out<=252;
				end
				if(in == 236) begin
					state<=17;
					out<=253;
				end
				if(in == 237) begin
					state<=1;
					out<=254;
				end
				if(in == 238) begin
					state<=17;
					out<=255;
				end
				if(in == 239) begin
					state<=17;
					out<=0;
				end
				if(in == 240) begin
					state<=17;
					out<=1;
				end
				if(in == 241) begin
					state<=17;
					out<=2;
				end
				if(in == 242) begin
					state<=17;
					out<=3;
				end
				if(in == 243) begin
					state<=17;
					out<=4;
				end
				if(in == 244) begin
					state<=17;
					out<=5;
				end
				if(in == 245) begin
					state<=17;
					out<=6;
				end
				if(in == 246) begin
					state<=17;
					out<=7;
				end
				if(in == 247) begin
					state<=17;
					out<=8;
				end
				if(in == 248) begin
					state<=17;
					out<=9;
				end
				if(in == 249) begin
					state<=17;
					out<=10;
				end
				if(in == 250) begin
					state<=17;
					out<=11;
				end
				if(in == 251) begin
					state<=17;
					out<=12;
				end
				if(in == 252) begin
					state<=17;
					out<=13;
				end
				if(in == 253) begin
					state<=17;
					out<=14;
				end
				if(in == 254) begin
					state<=17;
					out<=15;
				end
				if(in == 255) begin
					state<=17;
					out<=16;
				end
				if(in == 256) begin
					state<=17;
					out<=17;
				end
				if(in == 257) begin
					state<=17;
					out<=18;
				end
				if(in == 258) begin
					state<=17;
					out<=19;
				end
				if(in == 259) begin
					state<=17;
					out<=20;
				end
				if(in == 260) begin
					state<=17;
					out<=21;
				end
				if(in == 261) begin
					state<=17;
					out<=22;
				end
				if(in == 262) begin
					state<=17;
					out<=23;
				end
				if(in == 263) begin
					state<=17;
					out<=24;
				end
				if(in == 264) begin
					state<=17;
					out<=25;
				end
				if(in == 265) begin
					state<=17;
					out<=26;
				end
				if(in == 266) begin
					state<=17;
					out<=27;
				end
				if(in == 267) begin
					state<=17;
					out<=28;
				end
				if(in == 268) begin
					state<=17;
					out<=29;
				end
				if(in == 269) begin
					state<=17;
					out<=30;
				end
				if(in == 270) begin
					state<=17;
					out<=31;
				end
				if(in == 271) begin
					state<=17;
					out<=32;
				end
				if(in == 272) begin
					state<=17;
					out<=33;
				end
				if(in == 273) begin
					state<=17;
					out<=34;
				end
				if(in == 274) begin
					state<=17;
					out<=35;
				end
				if(in == 275) begin
					state<=17;
					out<=36;
				end
				if(in == 276) begin
					state<=17;
					out<=37;
				end
				if(in == 277) begin
					state<=17;
					out<=38;
				end
				if(in == 278) begin
					state<=17;
					out<=39;
				end
				if(in == 279) begin
					state<=17;
					out<=40;
				end
				if(in == 280) begin
					state<=17;
					out<=41;
				end
				if(in == 281) begin
					state<=17;
					out<=42;
				end
				if(in == 282) begin
					state<=17;
					out<=43;
				end
				if(in == 283) begin
					state<=17;
					out<=44;
				end
				if(in == 284) begin
					state<=17;
					out<=45;
				end
				if(in == 285) begin
					state<=1;
					out<=46;
				end
				if(in == 286) begin
					state<=17;
					out<=47;
				end
				if(in == 287) begin
					state<=1;
					out<=48;
				end
				if(in == 288) begin
					state<=17;
					out<=49;
				end
				if(in == 289) begin
					state<=1;
					out<=50;
				end
				if(in == 290) begin
					state<=17;
					out<=51;
				end
				if(in == 291) begin
					state<=17;
					out<=52;
				end
				if(in == 292) begin
					state<=17;
					out<=53;
				end
				if(in == 293) begin
					state<=17;
					out<=54;
				end
				if(in == 294) begin
					state<=17;
					out<=55;
				end
				if(in == 295) begin
					state<=17;
					out<=56;
				end
				if(in == 296) begin
					state<=17;
					out<=57;
				end
				if(in == 297) begin
					state<=17;
					out<=58;
				end
				if(in == 298) begin
					state<=17;
					out<=59;
				end
				if(in == 299) begin
					state<=17;
					out<=60;
				end
				if(in == 300) begin
					state<=17;
					out<=61;
				end
				if(in == 301) begin
					state<=17;
					out<=62;
				end
				if(in == 302) begin
					state<=17;
					out<=63;
				end
				if(in == 303) begin
					state<=17;
					out<=64;
				end
				if(in == 304) begin
					state<=17;
					out<=65;
				end
				if(in == 305) begin
					state<=17;
					out<=66;
				end
				if(in == 306) begin
					state<=17;
					out<=67;
				end
				if(in == 307) begin
					state<=17;
					out<=68;
				end
				if(in == 308) begin
					state<=17;
					out<=69;
				end
				if(in == 309) begin
					state<=17;
					out<=70;
				end
				if(in == 310) begin
					state<=17;
					out<=71;
				end
				if(in == 311) begin
					state<=17;
					out<=72;
				end
				if(in == 312) begin
					state<=17;
					out<=73;
				end
				if(in == 313) begin
					state<=17;
					out<=74;
				end
				if(in == 314) begin
					state<=17;
					out<=75;
				end
				if(in == 315) begin
					state<=17;
					out<=76;
				end
				if(in == 316) begin
					state<=17;
					out<=77;
				end
				if(in == 317) begin
					state<=17;
					out<=78;
				end
				if(in == 318) begin
					state<=17;
					out<=79;
				end
				if(in == 319) begin
					state<=17;
					out<=80;
				end
				if(in == 320) begin
					state<=17;
					out<=81;
				end
				if(in == 321) begin
					state<=17;
					out<=82;
				end
				if(in == 322) begin
					state<=17;
					out<=83;
				end
				if(in == 323) begin
					state<=17;
					out<=84;
				end
				if(in == 324) begin
					state<=17;
					out<=85;
				end
				if(in == 325) begin
					state<=17;
					out<=86;
				end
				if(in == 326) begin
					state<=17;
					out<=87;
				end
				if(in == 327) begin
					state<=17;
					out<=88;
				end
				if(in == 328) begin
					state<=17;
					out<=89;
				end
				if(in == 329) begin
					state<=17;
					out<=90;
				end
				if(in == 330) begin
					state<=17;
					out<=91;
				end
				if(in == 331) begin
					state<=17;
					out<=92;
				end
				if(in == 332) begin
					state<=17;
					out<=93;
				end
				if(in == 333) begin
					state<=17;
					out<=94;
				end
				if(in == 334) begin
					state<=17;
					out<=95;
				end
				if(in == 335) begin
					state<=17;
					out<=96;
				end
				if(in == 336) begin
					state<=17;
					out<=97;
				end
				if(in == 337) begin
					state<=1;
					out<=98;
				end
				if(in == 338) begin
					state<=17;
					out<=99;
				end
				if(in == 339) begin
					state<=1;
					out<=100;
				end
				if(in == 340) begin
					state<=17;
					out<=101;
				end
				if(in == 341) begin
					state<=1;
					out<=102;
				end
				if(in == 342) begin
					state<=17;
					out<=103;
				end
				if(in == 343) begin
					state<=1;
					out<=104;
				end
				if(in == 344) begin
					state<=17;
					out<=105;
				end
				if(in == 345) begin
					state<=1;
					out<=106;
				end
				if(in == 346) begin
					state<=17;
					out<=107;
				end
				if(in == 347) begin
					state<=1;
					out<=108;
				end
				if(in == 348) begin
					state<=17;
					out<=109;
				end
				if(in == 349) begin
					state<=1;
					out<=110;
				end
				if(in == 350) begin
					state<=17;
					out<=111;
				end
				if(in == 351) begin
					state<=1;
					out<=112;
				end
				if(in == 352) begin
					state<=17;
					out<=113;
				end
				if(in == 353) begin
					state<=1;
					out<=114;
				end
				if(in == 354) begin
					state<=17;
					out<=115;
				end
				if(in == 355) begin
					state<=17;
					out<=116;
				end
				if(in == 356) begin
					state<=17;
					out<=117;
				end
				if(in == 357) begin
					state<=17;
					out<=118;
				end
				if(in == 358) begin
					state<=17;
					out<=119;
				end
				if(in == 359) begin
					state<=17;
					out<=120;
				end
				if(in == 360) begin
					state<=17;
					out<=121;
				end
				if(in == 361) begin
					state<=17;
					out<=122;
				end
				if(in == 362) begin
					state<=17;
					out<=123;
				end
				if(in == 363) begin
					state<=17;
					out<=124;
				end
				if(in == 364) begin
					state<=17;
					out<=125;
				end
				if(in == 365) begin
					state<=17;
					out<=126;
				end
				if(in == 366) begin
					state<=17;
					out<=127;
				end
				if(in == 367) begin
					state<=17;
					out<=128;
				end
				if(in == 368) begin
					state<=17;
					out<=129;
				end
				if(in == 369) begin
					state<=17;
					out<=130;
				end
				if(in == 370) begin
					state<=17;
					out<=131;
				end
				if(in == 371) begin
					state<=17;
					out<=132;
				end
				if(in == 372) begin
					state<=17;
					out<=133;
				end
				if(in == 373) begin
					state<=17;
					out<=134;
				end
				if(in == 374) begin
					state<=17;
					out<=135;
				end
				if(in == 375) begin
					state<=17;
					out<=136;
				end
				if(in == 376) begin
					state<=17;
					out<=137;
				end
				if(in == 377) begin
					state<=17;
					out<=138;
				end
				if(in == 378) begin
					state<=17;
					out<=139;
				end
				if(in == 379) begin
					state<=17;
					out<=140;
				end
				if(in == 380) begin
					state<=17;
					out<=141;
				end
				if(in == 381) begin
					state<=17;
					out<=142;
				end
				if(in == 382) begin
					state<=17;
					out<=143;
				end
				if(in == 383) begin
					state<=17;
					out<=144;
				end
				if(in == 384) begin
					state<=17;
					out<=145;
				end
				if(in == 385) begin
					state<=17;
					out<=146;
				end
				if(in == 386) begin
					state<=17;
					out<=147;
				end
				if(in == 387) begin
					state<=17;
					out<=148;
				end
				if(in == 388) begin
					state<=17;
					out<=149;
				end
				if(in == 389) begin
					state<=17;
					out<=150;
				end
				if(in == 390) begin
					state<=17;
					out<=151;
				end
				if(in == 391) begin
					state<=17;
					out<=152;
				end
				if(in == 392) begin
					state<=17;
					out<=153;
				end
				if(in == 393) begin
					state<=17;
					out<=154;
				end
				if(in == 394) begin
					state<=17;
					out<=155;
				end
				if(in == 395) begin
					state<=17;
					out<=156;
				end
				if(in == 396) begin
					state<=17;
					out<=157;
				end
				if(in == 397) begin
					state<=17;
					out<=158;
				end
				if(in == 398) begin
					state<=17;
					out<=159;
				end
				if(in == 399) begin
					state<=17;
					out<=160;
				end
				if(in == 400) begin
					state<=17;
					out<=161;
				end
				if(in == 401) begin
					state<=1;
					out<=162;
				end
				if(in == 402) begin
					state<=17;
					out<=163;
				end
				if(in == 403) begin
					state<=1;
					out<=164;
				end
				if(in == 404) begin
					state<=17;
					out<=165;
				end
				if(in == 405) begin
					state<=1;
					out<=166;
				end
				if(in == 406) begin
					state<=17;
					out<=167;
				end
				if(in == 407) begin
					state<=17;
					out<=168;
				end
				if(in == 408) begin
					state<=17;
					out<=169;
				end
				if(in == 409) begin
					state<=17;
					out<=170;
				end
				if(in == 410) begin
					state<=17;
					out<=171;
				end
				if(in == 411) begin
					state<=17;
					out<=172;
				end
				if(in == 412) begin
					state<=17;
					out<=173;
				end
				if(in == 413) begin
					state<=17;
					out<=174;
				end
				if(in == 414) begin
					state<=17;
					out<=175;
				end
				if(in == 415) begin
					state<=17;
					out<=176;
				end
				if(in == 416) begin
					state<=17;
					out<=177;
				end
				if(in == 417) begin
					state<=17;
					out<=178;
				end
				if(in == 418) begin
					state<=17;
					out<=179;
				end
				if(in == 419) begin
					state<=17;
					out<=180;
				end
				if(in == 420) begin
					state<=17;
					out<=181;
				end
				if(in == 421) begin
					state<=17;
					out<=182;
				end
				if(in == 422) begin
					state<=17;
					out<=183;
				end
				if(in == 423) begin
					state<=17;
					out<=184;
				end
				if(in == 424) begin
					state<=17;
					out<=185;
				end
				if(in == 425) begin
					state<=17;
					out<=186;
				end
				if(in == 426) begin
					state<=17;
					out<=187;
				end
				if(in == 427) begin
					state<=17;
					out<=188;
				end
				if(in == 428) begin
					state<=17;
					out<=189;
				end
				if(in == 429) begin
					state<=17;
					out<=190;
				end
				if(in == 430) begin
					state<=17;
					out<=191;
				end
				if(in == 431) begin
					state<=17;
					out<=192;
				end
				if(in == 432) begin
					state<=17;
					out<=193;
				end
				if(in == 433) begin
					state<=17;
					out<=194;
				end
				if(in == 434) begin
					state<=17;
					out<=195;
				end
				if(in == 435) begin
					state<=17;
					out<=196;
				end
				if(in == 436) begin
					state<=17;
					out<=197;
				end
				if(in == 437) begin
					state<=17;
					out<=198;
				end
				if(in == 438) begin
					state<=17;
					out<=199;
				end
				if(in == 439) begin
					state<=17;
					out<=200;
				end
				if(in == 440) begin
					state<=17;
					out<=201;
				end
				if(in == 441) begin
					state<=17;
					out<=202;
				end
				if(in == 442) begin
					state<=17;
					out<=203;
				end
				if(in == 443) begin
					state<=17;
					out<=204;
				end
				if(in == 444) begin
					state<=17;
					out<=205;
				end
				if(in == 445) begin
					state<=17;
					out<=206;
				end
				if(in == 446) begin
					state<=17;
					out<=207;
				end
				if(in == 447) begin
					state<=17;
					out<=208;
				end
				if(in == 448) begin
					state<=17;
					out<=209;
				end
				if(in == 449) begin
					state<=17;
					out<=210;
				end
				if(in == 450) begin
					state<=17;
					out<=211;
				end
				if(in == 451) begin
					state<=17;
					out<=212;
				end
				if(in == 452) begin
					state<=17;
					out<=213;
				end
				if(in == 453) begin
					state<=1;
					out<=214;
				end
				if(in == 454) begin
					state<=17;
					out<=215;
				end
				if(in == 455) begin
					state<=1;
					out<=216;
				end
				if(in == 456) begin
					state<=17;
					out<=217;
				end
				if(in == 457) begin
					state<=1;
					out<=218;
				end
				if(in == 458) begin
					state<=17;
					out<=219;
				end
				if(in == 459) begin
					state<=1;
					out<=220;
				end
				if(in == 460) begin
					state<=17;
					out<=221;
				end
				if(in == 461) begin
					state<=1;
					out<=222;
				end
				if(in == 462) begin
					state<=17;
					out<=223;
				end
				if(in == 463) begin
					state<=1;
					out<=224;
				end
				if(in == 464) begin
					state<=17;
					out<=225;
				end
				if(in == 465) begin
					state<=1;
					out<=226;
				end
				if(in == 466) begin
					state<=17;
					out<=227;
				end
				if(in == 467) begin
					state<=1;
					out<=228;
				end
				if(in == 468) begin
					state<=17;
					out<=229;
				end
				if(in == 469) begin
					state<=1;
					out<=230;
				end
				if(in == 470) begin
					state<=17;
					out<=231;
				end
				if(in == 471) begin
					state<=17;
					out<=232;
				end
				if(in == 472) begin
					state<=17;
					out<=233;
				end
				if(in == 473) begin
					state<=17;
					out<=234;
				end
				if(in == 474) begin
					state<=17;
					out<=235;
				end
				if(in == 475) begin
					state<=17;
					out<=236;
				end
				if(in == 476) begin
					state<=17;
					out<=237;
				end
				if(in == 477) begin
					state<=17;
					out<=238;
				end
				if(in == 478) begin
					state<=17;
					out<=239;
				end
				if(in == 479) begin
					state<=17;
					out<=240;
				end
				if(in == 480) begin
					state<=17;
					out<=241;
				end
				if(in == 481) begin
					state<=17;
					out<=242;
				end
				if(in == 482) begin
					state<=17;
					out<=243;
				end
				if(in == 483) begin
					state<=17;
					out<=244;
				end
				if(in == 484) begin
					state<=17;
					out<=245;
				end
				if(in == 485) begin
					state<=17;
					out<=246;
				end
				if(in == 486) begin
					state<=17;
					out<=247;
				end
				if(in == 487) begin
					state<=17;
					out<=248;
				end
				if(in == 488) begin
					state<=17;
					out<=249;
				end
				if(in == 489) begin
					state<=17;
					out<=250;
				end
				if(in == 490) begin
					state<=17;
					out<=251;
				end
				if(in == 491) begin
					state<=17;
					out<=252;
				end
				if(in == 492) begin
					state<=17;
					out<=253;
				end
				if(in == 493) begin
					state<=17;
					out<=254;
				end
				if(in == 494) begin
					state<=17;
					out<=255;
				end
				if(in == 495) begin
					state<=17;
					out<=0;
				end
				if(in == 496) begin
					state<=17;
					out<=1;
				end
				if(in == 497) begin
					state<=17;
					out<=2;
				end
				if(in == 498) begin
					state<=17;
					out<=3;
				end
				if(in == 499) begin
					state<=17;
					out<=4;
				end
				if(in == 500) begin
					state<=17;
					out<=5;
				end
				if(in == 501) begin
					state<=17;
					out<=6;
				end
				if(in == 502) begin
					state<=17;
					out<=7;
				end
				if(in == 503) begin
					state<=17;
					out<=8;
				end
				if(in == 504) begin
					state<=17;
					out<=9;
				end
				if(in == 505) begin
					state<=17;
					out<=10;
				end
				if(in == 506) begin
					state<=17;
					out<=11;
				end
				if(in == 507) begin
					state<=17;
					out<=12;
				end
				if(in == 508) begin
					state<=17;
					out<=13;
				end
				if(in == 509) begin
					state<=17;
					out<=14;
				end
				if(in == 510) begin
					state<=17;
					out<=15;
				end
				if(in == 511) begin
					state<=17;
					out<=16;
				end
				if(in == 512) begin
					state<=17;
					out<=17;
				end
				if(in == 513) begin
					state<=17;
					out<=18;
				end
				if(in == 514) begin
					state<=17;
					out<=19;
				end
				if(in == 515) begin
					state<=17;
					out<=20;
				end
				if(in == 516) begin
					state<=17;
					out<=21;
				end
				if(in == 517) begin
					state<=1;
					out<=22;
				end
				if(in == 518) begin
					state<=17;
					out<=23;
				end
				if(in == 519) begin
					state<=1;
					out<=24;
				end
				if(in == 520) begin
					state<=17;
					out<=25;
				end
				if(in == 521) begin
					state<=1;
					out<=26;
				end
				if(in == 522) begin
					state<=17;
					out<=27;
				end
				if(in == 523) begin
					state<=17;
					out<=28;
				end
				if(in == 524) begin
					state<=17;
					out<=29;
				end
				if(in == 525) begin
					state<=17;
					out<=30;
				end
				if(in == 526) begin
					state<=17;
					out<=31;
				end
				if(in == 527) begin
					state<=17;
					out<=32;
				end
				if(in == 528) begin
					state<=17;
					out<=33;
				end
				if(in == 529) begin
					state<=17;
					out<=34;
				end
				if(in == 530) begin
					state<=17;
					out<=35;
				end
				if(in == 531) begin
					state<=17;
					out<=36;
				end
				if(in == 532) begin
					state<=17;
					out<=37;
				end
				if(in == 533) begin
					state<=17;
					out<=38;
				end
				if(in == 534) begin
					state<=17;
					out<=39;
				end
				if(in == 535) begin
					state<=17;
					out<=40;
				end
				if(in == 536) begin
					state<=17;
					out<=41;
				end
				if(in == 537) begin
					state<=17;
					out<=42;
				end
				if(in == 538) begin
					state<=17;
					out<=43;
				end
				if(in == 539) begin
					state<=17;
					out<=44;
				end
				if(in == 540) begin
					state<=17;
					out<=45;
				end
				if(in == 541) begin
					state<=17;
					out<=46;
				end
				if(in == 542) begin
					state<=17;
					out<=47;
				end
				if(in == 543) begin
					state<=17;
					out<=48;
				end
				if(in == 544) begin
					state<=17;
					out<=49;
				end
				if(in == 545) begin
					state<=17;
					out<=50;
				end
				if(in == 546) begin
					state<=17;
					out<=51;
				end
				if(in == 547) begin
					state<=17;
					out<=52;
				end
				if(in == 548) begin
					state<=17;
					out<=53;
				end
				if(in == 549) begin
					state<=17;
					out<=54;
				end
				if(in == 550) begin
					state<=17;
					out<=55;
				end
				if(in == 551) begin
					state<=17;
					out<=56;
				end
				if(in == 552) begin
					state<=17;
					out<=57;
				end
				if(in == 553) begin
					state<=17;
					out<=58;
				end
				if(in == 554) begin
					state<=17;
					out<=59;
				end
				if(in == 555) begin
					state<=17;
					out<=60;
				end
				if(in == 556) begin
					state<=17;
					out<=61;
				end
				if(in == 557) begin
					state<=17;
					out<=62;
				end
				if(in == 558) begin
					state<=17;
					out<=63;
				end
				if(in == 559) begin
					state<=17;
					out<=64;
				end
				if(in == 560) begin
					state<=17;
					out<=65;
				end
				if(in == 561) begin
					state<=17;
					out<=66;
				end
				if(in == 562) begin
					state<=17;
					out<=67;
				end
				if(in == 563) begin
					state<=17;
					out<=68;
				end
				if(in == 564) begin
					state<=17;
					out<=69;
				end
				if(in == 565) begin
					state<=17;
					out<=70;
				end
				if(in == 566) begin
					state<=17;
					out<=71;
				end
				if(in == 567) begin
					state<=17;
					out<=72;
				end
				if(in == 568) begin
					state<=17;
					out<=73;
				end
				if(in == 569) begin
					state<=1;
					out<=74;
				end
				if(in == 570) begin
					state<=17;
					out<=75;
				end
				if(in == 571) begin
					state<=1;
					out<=76;
				end
				if(in == 572) begin
					state<=17;
					out<=77;
				end
				if(in == 573) begin
					state<=1;
					out<=78;
				end
				if(in == 574) begin
					state<=17;
					out<=79;
				end
				if(in == 575) begin
					state<=1;
					out<=80;
				end
				if(in == 576) begin
					state<=17;
					out<=81;
				end
				if(in == 577) begin
					state<=1;
					out<=82;
				end
				if(in == 578) begin
					state<=17;
					out<=83;
				end
				if(in == 579) begin
					state<=1;
					out<=84;
				end
				if(in == 580) begin
					state<=17;
					out<=85;
				end
				if(in == 581) begin
					state<=1;
					out<=86;
				end
				if(in == 582) begin
					state<=17;
					out<=87;
				end
				if(in == 583) begin
					state<=1;
					out<=88;
				end
				if(in == 584) begin
					state<=17;
					out<=89;
				end
				if(in == 585) begin
					state<=1;
					out<=90;
				end
				if(in == 586) begin
					state<=17;
					out<=91;
				end
				if(in == 587) begin
					state<=17;
					out<=92;
				end
				if(in == 588) begin
					state<=17;
					out<=93;
				end
				if(in == 589) begin
					state<=17;
					out<=94;
				end
				if(in == 590) begin
					state<=17;
					out<=95;
				end
				if(in == 591) begin
					state<=17;
					out<=96;
				end
				if(in == 592) begin
					state<=17;
					out<=97;
				end
				if(in == 593) begin
					state<=17;
					out<=98;
				end
				if(in == 594) begin
					state<=17;
					out<=99;
				end
				if(in == 595) begin
					state<=17;
					out<=100;
				end
				if(in == 596) begin
					state<=17;
					out<=101;
				end
				if(in == 597) begin
					state<=17;
					out<=102;
				end
				if(in == 598) begin
					state<=17;
					out<=103;
				end
				if(in == 599) begin
					state<=17;
					out<=104;
				end
				if(in == 600) begin
					state<=17;
					out<=105;
				end
				if(in == 601) begin
					state<=17;
					out<=106;
				end
				if(in == 602) begin
					state<=17;
					out<=107;
				end
				if(in == 603) begin
					state<=17;
					out<=108;
				end
				if(in == 604) begin
					state<=17;
					out<=109;
				end
				if(in == 605) begin
					state<=17;
					out<=110;
				end
				if(in == 606) begin
					state<=17;
					out<=111;
				end
				if(in == 607) begin
					state<=17;
					out<=112;
				end
				if(in == 608) begin
					state<=17;
					out<=113;
				end
				if(in == 609) begin
					state<=17;
					out<=114;
				end
				if(in == 610) begin
					state<=17;
					out<=115;
				end
				if(in == 611) begin
					state<=17;
					out<=116;
				end
				if(in == 612) begin
					state<=17;
					out<=117;
				end
				if(in == 613) begin
					state<=17;
					out<=118;
				end
				if(in == 614) begin
					state<=17;
					out<=119;
				end
				if(in == 615) begin
					state<=17;
					out<=120;
				end
				if(in == 616) begin
					state<=17;
					out<=121;
				end
				if(in == 617) begin
					state<=17;
					out<=122;
				end
				if(in == 618) begin
					state<=17;
					out<=123;
				end
				if(in == 619) begin
					state<=17;
					out<=124;
				end
				if(in == 620) begin
					state<=17;
					out<=125;
				end
				if(in == 621) begin
					state<=17;
					out<=126;
				end
				if(in == 622) begin
					state<=17;
					out<=127;
				end
				if(in == 623) begin
					state<=17;
					out<=128;
				end
				if(in == 624) begin
					state<=17;
					out<=129;
				end
				if(in == 625) begin
					state<=17;
					out<=130;
				end
				if(in == 626) begin
					state<=17;
					out<=131;
				end
				if(in == 627) begin
					state<=17;
					out<=132;
				end
				if(in == 628) begin
					state<=17;
					out<=133;
				end
				if(in == 629) begin
					state<=17;
					out<=134;
				end
				if(in == 630) begin
					state<=17;
					out<=135;
				end
				if(in == 631) begin
					state<=17;
					out<=136;
				end
				if(in == 632) begin
					state<=17;
					out<=137;
				end
				if(in == 633) begin
					state<=1;
					out<=138;
				end
				if(in == 634) begin
					state<=17;
					out<=139;
				end
				if(in == 635) begin
					state<=1;
					out<=140;
				end
				if(in == 636) begin
					state<=17;
					out<=141;
				end
				if(in == 637) begin
					state<=1;
					out<=142;
				end
				if(in == 638) begin
					state<=17;
					out<=143;
				end
				if(in == 639) begin
					state<=17;
					out<=144;
				end
				if(in == 640) begin
					state<=17;
					out<=145;
				end
				if(in == 641) begin
					state<=17;
					out<=146;
				end
				if(in == 642) begin
					state<=17;
					out<=147;
				end
				if(in == 643) begin
					state<=17;
					out<=148;
				end
				if(in == 644) begin
					state<=17;
					out<=149;
				end
				if(in == 645) begin
					state<=17;
					out<=150;
				end
				if(in == 646) begin
					state<=17;
					out<=151;
				end
				if(in == 647) begin
					state<=17;
					out<=152;
				end
				if(in == 648) begin
					state<=17;
					out<=153;
				end
				if(in == 649) begin
					state<=17;
					out<=154;
				end
				if(in == 650) begin
					state<=17;
					out<=155;
				end
				if(in == 651) begin
					state<=17;
					out<=156;
				end
				if(in == 652) begin
					state<=17;
					out<=157;
				end
				if(in == 653) begin
					state<=17;
					out<=158;
				end
				if(in == 654) begin
					state<=17;
					out<=159;
				end
				if(in == 655) begin
					state<=17;
					out<=160;
				end
				if(in == 656) begin
					state<=17;
					out<=161;
				end
				if(in == 657) begin
					state<=17;
					out<=162;
				end
				if(in == 658) begin
					state<=17;
					out<=163;
				end
				if(in == 659) begin
					state<=17;
					out<=164;
				end
				if(in == 660) begin
					state<=17;
					out<=165;
				end
				if(in == 661) begin
					state<=17;
					out<=166;
				end
				if(in == 662) begin
					state<=17;
					out<=167;
				end
				if(in == 663) begin
					state<=17;
					out<=168;
				end
				if(in == 664) begin
					state<=17;
					out<=169;
				end
				if(in == 665) begin
					state<=17;
					out<=170;
				end
				if(in == 666) begin
					state<=17;
					out<=171;
				end
				if(in == 667) begin
					state<=17;
					out<=172;
				end
				if(in == 668) begin
					state<=17;
					out<=173;
				end
				if(in == 669) begin
					state<=17;
					out<=174;
				end
				if(in == 670) begin
					state<=17;
					out<=175;
				end
				if(in == 671) begin
					state<=17;
					out<=176;
				end
				if(in == 672) begin
					state<=17;
					out<=177;
				end
				if(in == 673) begin
					state<=17;
					out<=178;
				end
				if(in == 674) begin
					state<=17;
					out<=179;
				end
				if(in == 675) begin
					state<=17;
					out<=180;
				end
				if(in == 676) begin
					state<=17;
					out<=181;
				end
				if(in == 677) begin
					state<=17;
					out<=182;
				end
				if(in == 678) begin
					state<=17;
					out<=183;
				end
				if(in == 679) begin
					state<=17;
					out<=184;
				end
				if(in == 680) begin
					state<=17;
					out<=185;
				end
				if(in == 681) begin
					state<=17;
					out<=186;
				end
				if(in == 682) begin
					state<=17;
					out<=187;
				end
				if(in == 683) begin
					state<=17;
					out<=188;
				end
				if(in == 684) begin
					state<=17;
					out<=189;
				end
				if(in == 685) begin
					state<=1;
					out<=190;
				end
				if(in == 686) begin
					state<=17;
					out<=191;
				end
				if(in == 687) begin
					state<=1;
					out<=192;
				end
				if(in == 688) begin
					state<=17;
					out<=193;
				end
				if(in == 689) begin
					state<=1;
					out<=194;
				end
				if(in == 690) begin
					state<=17;
					out<=195;
				end
				if(in == 691) begin
					state<=1;
					out<=196;
				end
				if(in == 692) begin
					state<=17;
					out<=197;
				end
				if(in == 693) begin
					state<=1;
					out<=198;
				end
				if(in == 694) begin
					state<=17;
					out<=199;
				end
				if(in == 695) begin
					state<=1;
					out<=200;
				end
				if(in == 696) begin
					state<=17;
					out<=201;
				end
				if(in == 697) begin
					state<=1;
					out<=202;
				end
				if(in == 698) begin
					state<=17;
					out<=203;
				end
				if(in == 699) begin
					state<=1;
					out<=204;
				end
				if(in == 700) begin
					state<=17;
					out<=205;
				end
				if(in == 701) begin
					state<=1;
					out<=206;
				end
				if(in == 702) begin
					state<=17;
					out<=207;
				end
				if(in == 703) begin
					state<=17;
					out<=208;
				end
				if(in == 704) begin
					state<=17;
					out<=209;
				end
				if(in == 705) begin
					state<=17;
					out<=210;
				end
				if(in == 706) begin
					state<=17;
					out<=211;
				end
				if(in == 707) begin
					state<=17;
					out<=212;
				end
				if(in == 708) begin
					state<=17;
					out<=213;
				end
				if(in == 709) begin
					state<=17;
					out<=214;
				end
				if(in == 710) begin
					state<=17;
					out<=215;
				end
				if(in == 711) begin
					state<=17;
					out<=216;
				end
				if(in == 712) begin
					state<=17;
					out<=217;
				end
				if(in == 713) begin
					state<=17;
					out<=218;
				end
				if(in == 714) begin
					state<=17;
					out<=219;
				end
				if(in == 715) begin
					state<=17;
					out<=220;
				end
				if(in == 716) begin
					state<=17;
					out<=221;
				end
				if(in == 717) begin
					state<=17;
					out<=222;
				end
				if(in == 718) begin
					state<=17;
					out<=223;
				end
				if(in == 719) begin
					state<=17;
					out<=224;
				end
				if(in == 720) begin
					state<=17;
					out<=225;
				end
				if(in == 721) begin
					state<=17;
					out<=226;
				end
				if(in == 722) begin
					state<=17;
					out<=227;
				end
				if(in == 723) begin
					state<=17;
					out<=228;
				end
				if(in == 724) begin
					state<=17;
					out<=229;
				end
				if(in == 725) begin
					state<=17;
					out<=230;
				end
				if(in == 726) begin
					state<=17;
					out<=231;
				end
				if(in == 727) begin
					state<=17;
					out<=232;
				end
				if(in == 728) begin
					state<=17;
					out<=233;
				end
				if(in == 729) begin
					state<=17;
					out<=234;
				end
				if(in == 730) begin
					state<=17;
					out<=235;
				end
				if(in == 731) begin
					state<=17;
					out<=236;
				end
				if(in == 732) begin
					state<=17;
					out<=237;
				end
				if(in == 733) begin
					state<=17;
					out<=238;
				end
				if(in == 734) begin
					state<=17;
					out<=239;
				end
				if(in == 735) begin
					state<=17;
					out<=240;
				end
				if(in == 736) begin
					state<=17;
					out<=241;
				end
				if(in == 737) begin
					state<=17;
					out<=242;
				end
				if(in == 738) begin
					state<=17;
					out<=243;
				end
				if(in == 739) begin
					state<=17;
					out<=244;
				end
				if(in == 740) begin
					state<=17;
					out<=245;
				end
				if(in == 741) begin
					state<=17;
					out<=246;
				end
				if(in == 742) begin
					state<=17;
					out<=247;
				end
				if(in == 743) begin
					state<=17;
					out<=248;
				end
				if(in == 744) begin
					state<=17;
					out<=249;
				end
				if(in == 745) begin
					state<=17;
					out<=250;
				end
				if(in == 746) begin
					state<=17;
					out<=251;
				end
				if(in == 747) begin
					state<=17;
					out<=252;
				end
				if(in == 748) begin
					state<=17;
					out<=253;
				end
				if(in == 749) begin
					state<=1;
					out<=254;
				end
				if(in == 750) begin
					state<=17;
					out<=255;
				end
				if(in == 751) begin
					state<=1;
					out<=0;
				end
				if(in == 752) begin
					state<=17;
					out<=1;
				end
				if(in == 753) begin
					state<=1;
					out<=2;
				end
				if(in == 754) begin
					state<=17;
					out<=3;
				end
				if(in == 755) begin
					state<=17;
					out<=4;
				end
				if(in == 756) begin
					state<=17;
					out<=5;
				end
				if(in == 757) begin
					state<=17;
					out<=6;
				end
				if(in == 758) begin
					state<=17;
					out<=7;
				end
				if(in == 759) begin
					state<=17;
					out<=8;
				end
				if(in == 760) begin
					state<=17;
					out<=9;
				end
				if(in == 761) begin
					state<=17;
					out<=10;
				end
				if(in == 762) begin
					state<=17;
					out<=11;
				end
				if(in == 763) begin
					state<=17;
					out<=12;
				end
				if(in == 764) begin
					state<=17;
					out<=13;
				end
				if(in == 765) begin
					state<=17;
					out<=14;
				end
				if(in == 766) begin
					state<=17;
					out<=15;
				end
				if(in == 767) begin
					state<=17;
					out<=16;
				end
				if(in == 768) begin
					state<=17;
					out<=17;
				end
				if(in == 769) begin
					state<=17;
					out<=18;
				end
				if(in == 770) begin
					state<=17;
					out<=19;
				end
				if(in == 771) begin
					state<=17;
					out<=20;
				end
				if(in == 772) begin
					state<=17;
					out<=21;
				end
				if(in == 773) begin
					state<=17;
					out<=22;
				end
				if(in == 774) begin
					state<=17;
					out<=23;
				end
				if(in == 775) begin
					state<=17;
					out<=24;
				end
				if(in == 776) begin
					state<=17;
					out<=25;
				end
				if(in == 777) begin
					state<=17;
					out<=26;
				end
				if(in == 778) begin
					state<=17;
					out<=27;
				end
				if(in == 779) begin
					state<=17;
					out<=28;
				end
				if(in == 780) begin
					state<=17;
					out<=29;
				end
				if(in == 781) begin
					state<=17;
					out<=30;
				end
				if(in == 782) begin
					state<=17;
					out<=31;
				end
				if(in == 783) begin
					state<=17;
					out<=32;
				end
				if(in == 784) begin
					state<=17;
					out<=33;
				end
				if(in == 785) begin
					state<=17;
					out<=34;
				end
				if(in == 786) begin
					state<=17;
					out<=35;
				end
				if(in == 787) begin
					state<=17;
					out<=36;
				end
				if(in == 788) begin
					state<=17;
					out<=37;
				end
				if(in == 789) begin
					state<=17;
					out<=38;
				end
				if(in == 790) begin
					state<=17;
					out<=39;
				end
				if(in == 791) begin
					state<=17;
					out<=40;
				end
				if(in == 792) begin
					state<=17;
					out<=41;
				end
				if(in == 793) begin
					state<=17;
					out<=42;
				end
				if(in == 794) begin
					state<=17;
					out<=43;
				end
				if(in == 795) begin
					state<=17;
					out<=44;
				end
				if(in == 796) begin
					state<=17;
					out<=45;
				end
				if(in == 797) begin
					state<=17;
					out<=46;
				end
				if(in == 798) begin
					state<=17;
					out<=47;
				end
				if(in == 799) begin
					state<=17;
					out<=48;
				end
				if(in == 800) begin
					state<=17;
					out<=49;
				end
				if(in == 801) begin
					state<=1;
					out<=50;
				end
				if(in == 802) begin
					state<=17;
					out<=51;
				end
				if(in == 803) begin
					state<=1;
					out<=52;
				end
				if(in == 804) begin
					state<=17;
					out<=53;
				end
				if(in == 805) begin
					state<=1;
					out<=54;
				end
				if(in == 806) begin
					state<=17;
					out<=55;
				end
				if(in == 807) begin
					state<=1;
					out<=56;
				end
				if(in == 808) begin
					state<=17;
					out<=57;
				end
				if(in == 809) begin
					state<=1;
					out<=58;
				end
				if(in == 810) begin
					state<=17;
					out<=59;
				end
				if(in == 811) begin
					state<=1;
					out<=60;
				end
				if(in == 812) begin
					state<=17;
					out<=61;
				end
				if(in == 813) begin
					state<=1;
					out<=62;
				end
				if(in == 814) begin
					state<=17;
					out<=63;
				end
				if(in == 815) begin
					state<=1;
					out<=64;
				end
				if(in == 816) begin
					state<=17;
					out<=65;
				end
				if(in == 817) begin
					state<=1;
					out<=66;
				end
				if(in == 818) begin
					state<=17;
					out<=67;
				end
				if(in == 819) begin
					state<=17;
					out<=68;
				end
				if(in == 820) begin
					state<=17;
					out<=69;
				end
				if(in == 821) begin
					state<=17;
					out<=70;
				end
				if(in == 822) begin
					state<=17;
					out<=71;
				end
				if(in == 823) begin
					state<=17;
					out<=72;
				end
				if(in == 824) begin
					state<=17;
					out<=73;
				end
				if(in == 825) begin
					state<=17;
					out<=74;
				end
				if(in == 826) begin
					state<=17;
					out<=75;
				end
				if(in == 827) begin
					state<=17;
					out<=76;
				end
				if(in == 828) begin
					state<=17;
					out<=77;
				end
				if(in == 829) begin
					state<=17;
					out<=78;
				end
				if(in == 830) begin
					state<=17;
					out<=79;
				end
				if(in == 831) begin
					state<=17;
					out<=80;
				end
				if(in == 832) begin
					state<=17;
					out<=81;
				end
				if(in == 833) begin
					state<=17;
					out<=82;
				end
				if(in == 834) begin
					state<=17;
					out<=83;
				end
				if(in == 835) begin
					state<=17;
					out<=84;
				end
				if(in == 836) begin
					state<=17;
					out<=85;
				end
				if(in == 837) begin
					state<=17;
					out<=86;
				end
				if(in == 838) begin
					state<=17;
					out<=87;
				end
				if(in == 839) begin
					state<=17;
					out<=88;
				end
				if(in == 840) begin
					state<=17;
					out<=89;
				end
				if(in == 841) begin
					state<=17;
					out<=90;
				end
				if(in == 842) begin
					state<=17;
					out<=91;
				end
				if(in == 843) begin
					state<=17;
					out<=92;
				end
				if(in == 844) begin
					state<=17;
					out<=93;
				end
				if(in == 845) begin
					state<=17;
					out<=94;
				end
				if(in == 846) begin
					state<=17;
					out<=95;
				end
				if(in == 847) begin
					state<=17;
					out<=96;
				end
				if(in == 848) begin
					state<=17;
					out<=97;
				end
				if(in == 849) begin
					state<=17;
					out<=98;
				end
				if(in == 850) begin
					state<=17;
					out<=99;
				end
				if(in == 851) begin
					state<=17;
					out<=100;
				end
				if(in == 852) begin
					state<=17;
					out<=101;
				end
				if(in == 853) begin
					state<=17;
					out<=102;
				end
				if(in == 854) begin
					state<=17;
					out<=103;
				end
				if(in == 855) begin
					state<=17;
					out<=104;
				end
				if(in == 856) begin
					state<=17;
					out<=105;
				end
				if(in == 857) begin
					state<=17;
					out<=106;
				end
				if(in == 858) begin
					state<=17;
					out<=107;
				end
				if(in == 859) begin
					state<=17;
					out<=108;
				end
				if(in == 860) begin
					state<=17;
					out<=109;
				end
				if(in == 861) begin
					state<=17;
					out<=110;
				end
				if(in == 862) begin
					state<=17;
					out<=111;
				end
				if(in == 863) begin
					state<=17;
					out<=112;
				end
				if(in == 864) begin
					state<=17;
					out<=113;
				end
				if(in == 865) begin
					state<=1;
					out<=114;
				end
				if(in == 866) begin
					state<=17;
					out<=115;
				end
				if(in == 867) begin
					state<=1;
					out<=116;
				end
				if(in == 868) begin
					state<=17;
					out<=117;
				end
				if(in == 869) begin
					state<=1;
					out<=118;
				end
				if(in == 870) begin
					state<=17;
					out<=119;
				end
				if(in == 871) begin
					state<=17;
					out<=120;
				end
				if(in == 872) begin
					state<=17;
					out<=121;
				end
				if(in == 873) begin
					state<=17;
					out<=122;
				end
				if(in == 874) begin
					state<=17;
					out<=123;
				end
				if(in == 875) begin
					state<=17;
					out<=124;
				end
				if(in == 876) begin
					state<=17;
					out<=125;
				end
				if(in == 877) begin
					state<=17;
					out<=126;
				end
				if(in == 878) begin
					state<=17;
					out<=127;
				end
				if(in == 879) begin
					state<=17;
					out<=128;
				end
				if(in == 880) begin
					state<=17;
					out<=129;
				end
				if(in == 881) begin
					state<=17;
					out<=130;
				end
				if(in == 882) begin
					state<=17;
					out<=131;
				end
				if(in == 883) begin
					state<=17;
					out<=132;
				end
				if(in == 884) begin
					state<=17;
					out<=133;
				end
				if(in == 885) begin
					state<=17;
					out<=134;
				end
				if(in == 886) begin
					state<=17;
					out<=135;
				end
				if(in == 887) begin
					state<=17;
					out<=136;
				end
				if(in == 888) begin
					state<=17;
					out<=137;
				end
				if(in == 889) begin
					state<=17;
					out<=138;
				end
				if(in == 890) begin
					state<=17;
					out<=139;
				end
				if(in == 891) begin
					state<=17;
					out<=140;
				end
				if(in == 892) begin
					state<=17;
					out<=141;
				end
				if(in == 893) begin
					state<=17;
					out<=142;
				end
				if(in == 894) begin
					state<=17;
					out<=143;
				end
				if(in == 895) begin
					state<=17;
					out<=144;
				end
				if(in == 896) begin
					state<=17;
					out<=145;
				end
				if(in == 897) begin
					state<=17;
					out<=146;
				end
				if(in == 898) begin
					state<=17;
					out<=147;
				end
				if(in == 899) begin
					state<=17;
					out<=148;
				end
				if(in == 900) begin
					state<=17;
					out<=149;
				end
				if(in == 901) begin
					state<=17;
					out<=150;
				end
				if(in == 902) begin
					state<=17;
					out<=151;
				end
				if(in == 903) begin
					state<=17;
					out<=152;
				end
				if(in == 904) begin
					state<=17;
					out<=153;
				end
				if(in == 905) begin
					state<=17;
					out<=154;
				end
				if(in == 906) begin
					state<=17;
					out<=155;
				end
				if(in == 907) begin
					state<=17;
					out<=156;
				end
				if(in == 908) begin
					state<=17;
					out<=157;
				end
				if(in == 909) begin
					state<=17;
					out<=158;
				end
				if(in == 910) begin
					state<=17;
					out<=159;
				end
				if(in == 911) begin
					state<=17;
					out<=160;
				end
				if(in == 912) begin
					state<=17;
					out<=161;
				end
				if(in == 913) begin
					state<=17;
					out<=162;
				end
				if(in == 914) begin
					state<=17;
					out<=163;
				end
				if(in == 915) begin
					state<=17;
					out<=164;
				end
				if(in == 916) begin
					state<=17;
					out<=165;
				end
				if(in == 917) begin
					state<=1;
					out<=166;
				end
				if(in == 918) begin
					state<=17;
					out<=167;
				end
				if(in == 919) begin
					state<=1;
					out<=168;
				end
				if(in == 920) begin
					state<=17;
					out<=169;
				end
				if(in == 921) begin
					state<=1;
					out<=170;
				end
				if(in == 922) begin
					state<=17;
					out<=171;
				end
				if(in == 923) begin
					state<=1;
					out<=172;
				end
				if(in == 924) begin
					state<=17;
					out<=173;
				end
				if(in == 925) begin
					state<=1;
					out<=174;
				end
				if(in == 926) begin
					state<=17;
					out<=175;
				end
				if(in == 927) begin
					state<=1;
					out<=176;
				end
				if(in == 928) begin
					state<=17;
					out<=177;
				end
			end
			18: begin
				if(in == 0) begin
					state<=3;
					out<=178;
				end
				if(in == 1) begin
					state<=1;
					out<=179;
				end
				if(in == 2) begin
					state<=18;
					out<=180;
				end
				if(in == 3) begin
					state<=3;
					out<=181;
				end
				if(in == 4) begin
					state<=22;
					out<=182;
				end
				if(in == 5) begin
					state<=3;
					out<=183;
				end
				if(in == 6) begin
					state<=22;
					out<=184;
				end
				if(in == 7) begin
					state<=19;
					out<=185;
				end
				if(in == 8) begin
					state<=19;
					out<=186;
				end
				if(in == 9) begin
					state<=22;
					out<=187;
				end
				if(in == 10) begin
					state<=22;
					out<=188;
				end
				if(in == 11) begin
					state<=19;
					out<=189;
				end
				if(in == 12) begin
					state<=19;
					out<=190;
				end
				if(in == 13) begin
					state<=22;
					out<=191;
				end
				if(in == 14) begin
					state<=22;
					out<=192;
				end
				if(in == 15) begin
					state<=19;
					out<=193;
				end
				if(in == 16) begin
					state<=19;
					out<=194;
				end
				if(in == 17) begin
					state<=22;
					out<=195;
				end
				if(in == 18) begin
					state<=22;
					out<=196;
				end
				if(in == 19) begin
					state<=19;
					out<=197;
				end
				if(in == 20) begin
					state<=19;
					out<=198;
				end
				if(in == 21) begin
					state<=22;
					out<=199;
				end
				if(in == 22) begin
					state<=22;
					out<=200;
				end
				if(in == 23) begin
					state<=19;
					out<=201;
				end
				if(in == 24) begin
					state<=19;
					out<=202;
				end
				if(in == 25) begin
					state<=22;
					out<=203;
				end
				if(in == 26) begin
					state<=22;
					out<=204;
				end
				if(in == 27) begin
					state<=19;
					out<=205;
				end
				if(in == 28) begin
					state<=19;
					out<=206;
				end
				if(in == 29) begin
					state<=22;
					out<=207;
				end
				if(in == 30) begin
					state<=22;
					out<=208;
				end
				if(in == 31) begin
					state<=19;
					out<=209;
				end
				if(in == 32) begin
					state<=19;
					out<=210;
				end
				if(in == 33) begin
					state<=22;
					out<=211;
				end
				if(in == 34) begin
					state<=22;
					out<=212;
				end
				if(in == 35) begin
					state<=19;
					out<=213;
				end
				if(in == 36) begin
					state<=19;
					out<=214;
				end
				if(in == 37) begin
					state<=22;
					out<=215;
				end
				if(in == 38) begin
					state<=22;
					out<=216;
				end
				if(in == 39) begin
					state<=19;
					out<=217;
				end
				if(in == 40) begin
					state<=19;
					out<=218;
				end
				if(in == 41) begin
					state<=22;
					out<=219;
				end
				if(in == 42) begin
					state<=22;
					out<=220;
				end
				if(in == 43) begin
					state<=19;
					out<=221;
				end
				if(in == 44) begin
					state<=19;
					out<=222;
				end
				if(in == 45) begin
					state<=22;
					out<=223;
				end
				if(in == 46) begin
					state<=22;
					out<=224;
				end
				if(in == 47) begin
					state<=19;
					out<=225;
				end
				if(in == 48) begin
					state<=19;
					out<=226;
				end
				if(in == 49) begin
					state<=22;
					out<=227;
				end
				if(in == 50) begin
					state<=22;
					out<=228;
				end
				if(in == 51) begin
					state<=19;
					out<=229;
				end
				if(in == 52) begin
					state<=19;
					out<=230;
				end
				if(in == 53) begin
					state<=3;
					out<=231;
				end
				if(in == 54) begin
					state<=18;
					out<=232;
				end
				if(in == 55) begin
					state<=3;
					out<=233;
				end
				if(in == 56) begin
					state<=22;
					out<=234;
				end
				if(in == 57) begin
					state<=3;
					out<=235;
				end
				if(in == 58) begin
					state<=22;
					out<=236;
				end
				if(in == 59) begin
					state<=19;
					out<=237;
				end
				if(in == 60) begin
					state<=19;
					out<=238;
				end
				if(in == 61) begin
					state<=22;
					out<=239;
				end
				if(in == 62) begin
					state<=22;
					out<=240;
				end
				if(in == 63) begin
					state<=19;
					out<=241;
				end
				if(in == 64) begin
					state<=19;
					out<=242;
				end
				if(in == 65) begin
					state<=22;
					out<=243;
				end
				if(in == 66) begin
					state<=22;
					out<=244;
				end
				if(in == 67) begin
					state<=19;
					out<=245;
				end
				if(in == 68) begin
					state<=19;
					out<=246;
				end
				if(in == 69) begin
					state<=22;
					out<=247;
				end
				if(in == 70) begin
					state<=22;
					out<=248;
				end
				if(in == 71) begin
					state<=19;
					out<=249;
				end
				if(in == 72) begin
					state<=19;
					out<=250;
				end
				if(in == 73) begin
					state<=22;
					out<=251;
				end
				if(in == 74) begin
					state<=22;
					out<=252;
				end
				if(in == 75) begin
					state<=19;
					out<=253;
				end
				if(in == 76) begin
					state<=19;
					out<=254;
				end
				if(in == 77) begin
					state<=22;
					out<=255;
				end
				if(in == 78) begin
					state<=22;
					out<=0;
				end
				if(in == 79) begin
					state<=19;
					out<=1;
				end
				if(in == 80) begin
					state<=19;
					out<=2;
				end
				if(in == 81) begin
					state<=22;
					out<=3;
				end
				if(in == 82) begin
					state<=22;
					out<=4;
				end
				if(in == 83) begin
					state<=19;
					out<=5;
				end
				if(in == 84) begin
					state<=19;
					out<=6;
				end
				if(in == 85) begin
					state<=22;
					out<=7;
				end
				if(in == 86) begin
					state<=22;
					out<=8;
				end
				if(in == 87) begin
					state<=19;
					out<=9;
				end
				if(in == 88) begin
					state<=19;
					out<=10;
				end
				if(in == 89) begin
					state<=22;
					out<=11;
				end
				if(in == 90) begin
					state<=22;
					out<=12;
				end
				if(in == 91) begin
					state<=19;
					out<=13;
				end
				if(in == 92) begin
					state<=19;
					out<=14;
				end
				if(in == 93) begin
					state<=22;
					out<=15;
				end
				if(in == 94) begin
					state<=22;
					out<=16;
				end
				if(in == 95) begin
					state<=19;
					out<=17;
				end
				if(in == 96) begin
					state<=19;
					out<=18;
				end
				if(in == 97) begin
					state<=22;
					out<=19;
				end
				if(in == 98) begin
					state<=22;
					out<=20;
				end
				if(in == 99) begin
					state<=19;
					out<=21;
				end
				if(in == 100) begin
					state<=19;
					out<=22;
				end
				if(in == 101) begin
					state<=22;
					out<=23;
				end
				if(in == 102) begin
					state<=22;
					out<=24;
				end
				if(in == 103) begin
					state<=19;
					out<=25;
				end
				if(in == 104) begin
					state<=19;
					out<=26;
				end
				if(in == 105) begin
					state<=2;
					out<=27;
				end
				if(in == 106) begin
					state<=2;
					out<=28;
				end
				if(in == 107) begin
					state<=2;
					out<=29;
				end
				if(in == 108) begin
					state<=2;
					out<=30;
				end
				if(in == 109) begin
					state<=2;
					out<=31;
				end
				if(in == 110) begin
					state<=2;
					out<=32;
				end
				if(in == 111) begin
					state<=2;
					out<=33;
				end
				if(in == 112) begin
					state<=2;
					out<=34;
				end
				if(in == 113) begin
					state<=2;
					out<=35;
				end
				if(in == 114) begin
					state<=2;
					out<=36;
				end
				if(in == 115) begin
					state<=2;
					out<=37;
				end
				if(in == 116) begin
					state<=2;
					out<=38;
				end
				if(in == 117) begin
					state<=3;
					out<=39;
				end
				if(in == 118) begin
					state<=18;
					out<=40;
				end
				if(in == 119) begin
					state<=3;
					out<=41;
				end
				if(in == 120) begin
					state<=22;
					out<=42;
				end
				if(in == 121) begin
					state<=3;
					out<=43;
				end
				if(in == 122) begin
					state<=22;
					out<=44;
				end
				if(in == 123) begin
					state<=19;
					out<=45;
				end
				if(in == 124) begin
					state<=19;
					out<=46;
				end
				if(in == 125) begin
					state<=22;
					out<=47;
				end
				if(in == 126) begin
					state<=22;
					out<=48;
				end
				if(in == 127) begin
					state<=19;
					out<=49;
				end
				if(in == 128) begin
					state<=19;
					out<=50;
				end
				if(in == 129) begin
					state<=22;
					out<=51;
				end
				if(in == 130) begin
					state<=22;
					out<=52;
				end
				if(in == 131) begin
					state<=19;
					out<=53;
				end
				if(in == 132) begin
					state<=19;
					out<=54;
				end
				if(in == 133) begin
					state<=22;
					out<=55;
				end
				if(in == 134) begin
					state<=22;
					out<=56;
				end
				if(in == 135) begin
					state<=19;
					out<=57;
				end
				if(in == 136) begin
					state<=19;
					out<=58;
				end
				if(in == 137) begin
					state<=22;
					out<=59;
				end
				if(in == 138) begin
					state<=22;
					out<=60;
				end
				if(in == 139) begin
					state<=19;
					out<=61;
				end
				if(in == 140) begin
					state<=19;
					out<=62;
				end
				if(in == 141) begin
					state<=22;
					out<=63;
				end
				if(in == 142) begin
					state<=22;
					out<=64;
				end
				if(in == 143) begin
					state<=19;
					out<=65;
				end
				if(in == 144) begin
					state<=19;
					out<=66;
				end
				if(in == 145) begin
					state<=22;
					out<=67;
				end
				if(in == 146) begin
					state<=22;
					out<=68;
				end
				if(in == 147) begin
					state<=19;
					out<=69;
				end
				if(in == 148) begin
					state<=19;
					out<=70;
				end
				if(in == 149) begin
					state<=22;
					out<=71;
				end
				if(in == 150) begin
					state<=22;
					out<=72;
				end
				if(in == 151) begin
					state<=19;
					out<=73;
				end
				if(in == 152) begin
					state<=19;
					out<=74;
				end
				if(in == 153) begin
					state<=22;
					out<=75;
				end
				if(in == 154) begin
					state<=22;
					out<=76;
				end
				if(in == 155) begin
					state<=19;
					out<=77;
				end
				if(in == 156) begin
					state<=19;
					out<=78;
				end
				if(in == 157) begin
					state<=22;
					out<=79;
				end
				if(in == 158) begin
					state<=22;
					out<=80;
				end
				if(in == 159) begin
					state<=19;
					out<=81;
				end
				if(in == 160) begin
					state<=19;
					out<=82;
				end
				if(in == 161) begin
					state<=22;
					out<=83;
				end
				if(in == 162) begin
					state<=22;
					out<=84;
				end
				if(in == 163) begin
					state<=19;
					out<=85;
				end
				if(in == 164) begin
					state<=19;
					out<=86;
				end
				if(in == 165) begin
					state<=22;
					out<=87;
				end
				if(in == 166) begin
					state<=22;
					out<=88;
				end
				if(in == 167) begin
					state<=19;
					out<=89;
				end
				if(in == 168) begin
					state<=19;
					out<=90;
				end
				if(in == 169) begin
					state<=3;
					out<=91;
				end
				if(in == 170) begin
					state<=18;
					out<=92;
				end
				if(in == 171) begin
					state<=3;
					out<=93;
				end
				if(in == 172) begin
					state<=22;
					out<=94;
				end
				if(in == 173) begin
					state<=3;
					out<=95;
				end
				if(in == 174) begin
					state<=22;
					out<=96;
				end
				if(in == 175) begin
					state<=19;
					out<=97;
				end
				if(in == 176) begin
					state<=19;
					out<=98;
				end
				if(in == 177) begin
					state<=22;
					out<=99;
				end
				if(in == 178) begin
					state<=22;
					out<=100;
				end
				if(in == 179) begin
					state<=19;
					out<=101;
				end
				if(in == 180) begin
					state<=19;
					out<=102;
				end
				if(in == 181) begin
					state<=22;
					out<=103;
				end
				if(in == 182) begin
					state<=22;
					out<=104;
				end
				if(in == 183) begin
					state<=19;
					out<=105;
				end
				if(in == 184) begin
					state<=19;
					out<=106;
				end
				if(in == 185) begin
					state<=22;
					out<=107;
				end
				if(in == 186) begin
					state<=22;
					out<=108;
				end
				if(in == 187) begin
					state<=19;
					out<=109;
				end
				if(in == 188) begin
					state<=19;
					out<=110;
				end
				if(in == 189) begin
					state<=22;
					out<=111;
				end
				if(in == 190) begin
					state<=22;
					out<=112;
				end
				if(in == 191) begin
					state<=19;
					out<=113;
				end
				if(in == 192) begin
					state<=19;
					out<=114;
				end
				if(in == 193) begin
					state<=22;
					out<=115;
				end
				if(in == 194) begin
					state<=22;
					out<=116;
				end
				if(in == 195) begin
					state<=19;
					out<=117;
				end
				if(in == 196) begin
					state<=19;
					out<=118;
				end
				if(in == 197) begin
					state<=22;
					out<=119;
				end
				if(in == 198) begin
					state<=22;
					out<=120;
				end
				if(in == 199) begin
					state<=19;
					out<=121;
				end
				if(in == 200) begin
					state<=19;
					out<=122;
				end
				if(in == 201) begin
					state<=22;
					out<=123;
				end
				if(in == 202) begin
					state<=22;
					out<=124;
				end
				if(in == 203) begin
					state<=19;
					out<=125;
				end
				if(in == 204) begin
					state<=19;
					out<=126;
				end
				if(in == 205) begin
					state<=22;
					out<=127;
				end
				if(in == 206) begin
					state<=22;
					out<=128;
				end
				if(in == 207) begin
					state<=19;
					out<=129;
				end
				if(in == 208) begin
					state<=19;
					out<=130;
				end
				if(in == 209) begin
					state<=22;
					out<=131;
				end
				if(in == 210) begin
					state<=22;
					out<=132;
				end
				if(in == 211) begin
					state<=19;
					out<=133;
				end
				if(in == 212) begin
					state<=19;
					out<=134;
				end
				if(in == 213) begin
					state<=22;
					out<=135;
				end
				if(in == 214) begin
					state<=22;
					out<=136;
				end
				if(in == 215) begin
					state<=19;
					out<=137;
				end
				if(in == 216) begin
					state<=19;
					out<=138;
				end
				if(in == 217) begin
					state<=22;
					out<=139;
				end
				if(in == 218) begin
					state<=22;
					out<=140;
				end
				if(in == 219) begin
					state<=19;
					out<=141;
				end
				if(in == 220) begin
					state<=19;
					out<=142;
				end
				if(in == 221) begin
					state<=2;
					out<=143;
				end
				if(in == 222) begin
					state<=2;
					out<=144;
				end
				if(in == 223) begin
					state<=2;
					out<=145;
				end
				if(in == 224) begin
					state<=2;
					out<=146;
				end
				if(in == 225) begin
					state<=2;
					out<=147;
				end
				if(in == 226) begin
					state<=2;
					out<=148;
				end
				if(in == 227) begin
					state<=2;
					out<=149;
				end
				if(in == 228) begin
					state<=2;
					out<=150;
				end
				if(in == 229) begin
					state<=2;
					out<=151;
				end
				if(in == 230) begin
					state<=2;
					out<=152;
				end
				if(in == 231) begin
					state<=2;
					out<=153;
				end
				if(in == 232) begin
					state<=2;
					out<=154;
				end
				if(in == 233) begin
					state<=3;
					out<=155;
				end
				if(in == 234) begin
					state<=18;
					out<=156;
				end
				if(in == 235) begin
					state<=3;
					out<=157;
				end
				if(in == 236) begin
					state<=22;
					out<=158;
				end
				if(in == 237) begin
					state<=3;
					out<=159;
				end
				if(in == 238) begin
					state<=22;
					out<=160;
				end
				if(in == 239) begin
					state<=19;
					out<=161;
				end
				if(in == 240) begin
					state<=19;
					out<=162;
				end
				if(in == 241) begin
					state<=22;
					out<=163;
				end
				if(in == 242) begin
					state<=22;
					out<=164;
				end
				if(in == 243) begin
					state<=19;
					out<=165;
				end
				if(in == 244) begin
					state<=19;
					out<=166;
				end
				if(in == 245) begin
					state<=22;
					out<=167;
				end
				if(in == 246) begin
					state<=22;
					out<=168;
				end
				if(in == 247) begin
					state<=19;
					out<=169;
				end
				if(in == 248) begin
					state<=19;
					out<=170;
				end
				if(in == 249) begin
					state<=22;
					out<=171;
				end
				if(in == 250) begin
					state<=22;
					out<=172;
				end
				if(in == 251) begin
					state<=19;
					out<=173;
				end
				if(in == 252) begin
					state<=19;
					out<=174;
				end
				if(in == 253) begin
					state<=22;
					out<=175;
				end
				if(in == 254) begin
					state<=22;
					out<=176;
				end
				if(in == 255) begin
					state<=19;
					out<=177;
				end
				if(in == 256) begin
					state<=19;
					out<=178;
				end
				if(in == 257) begin
					state<=22;
					out<=179;
				end
				if(in == 258) begin
					state<=22;
					out<=180;
				end
				if(in == 259) begin
					state<=19;
					out<=181;
				end
				if(in == 260) begin
					state<=19;
					out<=182;
				end
				if(in == 261) begin
					state<=22;
					out<=183;
				end
				if(in == 262) begin
					state<=22;
					out<=184;
				end
				if(in == 263) begin
					state<=19;
					out<=185;
				end
				if(in == 264) begin
					state<=19;
					out<=186;
				end
				if(in == 265) begin
					state<=22;
					out<=187;
				end
				if(in == 266) begin
					state<=22;
					out<=188;
				end
				if(in == 267) begin
					state<=19;
					out<=189;
				end
				if(in == 268) begin
					state<=19;
					out<=190;
				end
				if(in == 269) begin
					state<=22;
					out<=191;
				end
				if(in == 270) begin
					state<=22;
					out<=192;
				end
				if(in == 271) begin
					state<=19;
					out<=193;
				end
				if(in == 272) begin
					state<=19;
					out<=194;
				end
				if(in == 273) begin
					state<=22;
					out<=195;
				end
				if(in == 274) begin
					state<=22;
					out<=196;
				end
				if(in == 275) begin
					state<=19;
					out<=197;
				end
				if(in == 276) begin
					state<=19;
					out<=198;
				end
				if(in == 277) begin
					state<=22;
					out<=199;
				end
				if(in == 278) begin
					state<=22;
					out<=200;
				end
				if(in == 279) begin
					state<=19;
					out<=201;
				end
				if(in == 280) begin
					state<=19;
					out<=202;
				end
				if(in == 281) begin
					state<=22;
					out<=203;
				end
				if(in == 282) begin
					state<=22;
					out<=204;
				end
				if(in == 283) begin
					state<=19;
					out<=205;
				end
				if(in == 284) begin
					state<=19;
					out<=206;
				end
				if(in == 285) begin
					state<=3;
					out<=207;
				end
				if(in == 286) begin
					state<=18;
					out<=208;
				end
				if(in == 287) begin
					state<=3;
					out<=209;
				end
				if(in == 288) begin
					state<=22;
					out<=210;
				end
				if(in == 289) begin
					state<=3;
					out<=211;
				end
				if(in == 290) begin
					state<=22;
					out<=212;
				end
				if(in == 291) begin
					state<=19;
					out<=213;
				end
				if(in == 292) begin
					state<=19;
					out<=214;
				end
				if(in == 293) begin
					state<=22;
					out<=215;
				end
				if(in == 294) begin
					state<=22;
					out<=216;
				end
				if(in == 295) begin
					state<=19;
					out<=217;
				end
				if(in == 296) begin
					state<=19;
					out<=218;
				end
				if(in == 297) begin
					state<=22;
					out<=219;
				end
				if(in == 298) begin
					state<=22;
					out<=220;
				end
				if(in == 299) begin
					state<=19;
					out<=221;
				end
				if(in == 300) begin
					state<=19;
					out<=222;
				end
				if(in == 301) begin
					state<=22;
					out<=223;
				end
				if(in == 302) begin
					state<=22;
					out<=224;
				end
				if(in == 303) begin
					state<=19;
					out<=225;
				end
				if(in == 304) begin
					state<=19;
					out<=226;
				end
				if(in == 305) begin
					state<=22;
					out<=227;
				end
				if(in == 306) begin
					state<=22;
					out<=228;
				end
				if(in == 307) begin
					state<=19;
					out<=229;
				end
				if(in == 308) begin
					state<=19;
					out<=230;
				end
				if(in == 309) begin
					state<=22;
					out<=231;
				end
				if(in == 310) begin
					state<=22;
					out<=232;
				end
				if(in == 311) begin
					state<=19;
					out<=233;
				end
				if(in == 312) begin
					state<=19;
					out<=234;
				end
				if(in == 313) begin
					state<=22;
					out<=235;
				end
				if(in == 314) begin
					state<=22;
					out<=236;
				end
				if(in == 315) begin
					state<=19;
					out<=237;
				end
				if(in == 316) begin
					state<=19;
					out<=238;
				end
				if(in == 317) begin
					state<=22;
					out<=239;
				end
				if(in == 318) begin
					state<=22;
					out<=240;
				end
				if(in == 319) begin
					state<=19;
					out<=241;
				end
				if(in == 320) begin
					state<=19;
					out<=242;
				end
				if(in == 321) begin
					state<=22;
					out<=243;
				end
				if(in == 322) begin
					state<=22;
					out<=244;
				end
				if(in == 323) begin
					state<=19;
					out<=245;
				end
				if(in == 324) begin
					state<=19;
					out<=246;
				end
				if(in == 325) begin
					state<=22;
					out<=247;
				end
				if(in == 326) begin
					state<=22;
					out<=248;
				end
				if(in == 327) begin
					state<=19;
					out<=249;
				end
				if(in == 328) begin
					state<=19;
					out<=250;
				end
				if(in == 329) begin
					state<=22;
					out<=251;
				end
				if(in == 330) begin
					state<=22;
					out<=252;
				end
				if(in == 331) begin
					state<=19;
					out<=253;
				end
				if(in == 332) begin
					state<=19;
					out<=254;
				end
				if(in == 333) begin
					state<=22;
					out<=255;
				end
				if(in == 334) begin
					state<=22;
					out<=0;
				end
				if(in == 335) begin
					state<=19;
					out<=1;
				end
				if(in == 336) begin
					state<=19;
					out<=2;
				end
				if(in == 337) begin
					state<=2;
					out<=3;
				end
				if(in == 338) begin
					state<=2;
					out<=4;
				end
				if(in == 339) begin
					state<=2;
					out<=5;
				end
				if(in == 340) begin
					state<=2;
					out<=6;
				end
				if(in == 341) begin
					state<=2;
					out<=7;
				end
				if(in == 342) begin
					state<=2;
					out<=8;
				end
				if(in == 343) begin
					state<=2;
					out<=9;
				end
				if(in == 344) begin
					state<=2;
					out<=10;
				end
				if(in == 345) begin
					state<=2;
					out<=11;
				end
				if(in == 346) begin
					state<=2;
					out<=12;
				end
				if(in == 347) begin
					state<=2;
					out<=13;
				end
				if(in == 348) begin
					state<=2;
					out<=14;
				end
				if(in == 349) begin
					state<=3;
					out<=15;
				end
				if(in == 350) begin
					state<=18;
					out<=16;
				end
				if(in == 351) begin
					state<=3;
					out<=17;
				end
				if(in == 352) begin
					state<=22;
					out<=18;
				end
				if(in == 353) begin
					state<=3;
					out<=19;
				end
				if(in == 354) begin
					state<=22;
					out<=20;
				end
				if(in == 355) begin
					state<=19;
					out<=21;
				end
				if(in == 356) begin
					state<=19;
					out<=22;
				end
				if(in == 357) begin
					state<=22;
					out<=23;
				end
				if(in == 358) begin
					state<=22;
					out<=24;
				end
				if(in == 359) begin
					state<=19;
					out<=25;
				end
				if(in == 360) begin
					state<=19;
					out<=26;
				end
				if(in == 361) begin
					state<=22;
					out<=27;
				end
				if(in == 362) begin
					state<=22;
					out<=28;
				end
				if(in == 363) begin
					state<=19;
					out<=29;
				end
				if(in == 364) begin
					state<=19;
					out<=30;
				end
				if(in == 365) begin
					state<=22;
					out<=31;
				end
				if(in == 366) begin
					state<=22;
					out<=32;
				end
				if(in == 367) begin
					state<=19;
					out<=33;
				end
				if(in == 368) begin
					state<=19;
					out<=34;
				end
				if(in == 369) begin
					state<=22;
					out<=35;
				end
				if(in == 370) begin
					state<=22;
					out<=36;
				end
				if(in == 371) begin
					state<=19;
					out<=37;
				end
				if(in == 372) begin
					state<=19;
					out<=38;
				end
				if(in == 373) begin
					state<=22;
					out<=39;
				end
				if(in == 374) begin
					state<=22;
					out<=40;
				end
				if(in == 375) begin
					state<=19;
					out<=41;
				end
				if(in == 376) begin
					state<=19;
					out<=42;
				end
				if(in == 377) begin
					state<=22;
					out<=43;
				end
				if(in == 378) begin
					state<=22;
					out<=44;
				end
				if(in == 379) begin
					state<=19;
					out<=45;
				end
				if(in == 380) begin
					state<=19;
					out<=46;
				end
				if(in == 381) begin
					state<=22;
					out<=47;
				end
				if(in == 382) begin
					state<=22;
					out<=48;
				end
				if(in == 383) begin
					state<=19;
					out<=49;
				end
				if(in == 384) begin
					state<=19;
					out<=50;
				end
				if(in == 385) begin
					state<=22;
					out<=51;
				end
				if(in == 386) begin
					state<=22;
					out<=52;
				end
				if(in == 387) begin
					state<=19;
					out<=53;
				end
				if(in == 388) begin
					state<=19;
					out<=54;
				end
				if(in == 389) begin
					state<=22;
					out<=55;
				end
				if(in == 390) begin
					state<=22;
					out<=56;
				end
				if(in == 391) begin
					state<=19;
					out<=57;
				end
				if(in == 392) begin
					state<=19;
					out<=58;
				end
				if(in == 393) begin
					state<=22;
					out<=59;
				end
				if(in == 394) begin
					state<=22;
					out<=60;
				end
				if(in == 395) begin
					state<=19;
					out<=61;
				end
				if(in == 396) begin
					state<=19;
					out<=62;
				end
				if(in == 397) begin
					state<=22;
					out<=63;
				end
				if(in == 398) begin
					state<=22;
					out<=64;
				end
				if(in == 399) begin
					state<=19;
					out<=65;
				end
				if(in == 400) begin
					state<=19;
					out<=66;
				end
				if(in == 401) begin
					state<=3;
					out<=67;
				end
				if(in == 402) begin
					state<=18;
					out<=68;
				end
				if(in == 403) begin
					state<=3;
					out<=69;
				end
				if(in == 404) begin
					state<=22;
					out<=70;
				end
				if(in == 405) begin
					state<=3;
					out<=71;
				end
				if(in == 406) begin
					state<=22;
					out<=72;
				end
				if(in == 407) begin
					state<=19;
					out<=73;
				end
				if(in == 408) begin
					state<=19;
					out<=74;
				end
				if(in == 409) begin
					state<=22;
					out<=75;
				end
				if(in == 410) begin
					state<=22;
					out<=76;
				end
				if(in == 411) begin
					state<=19;
					out<=77;
				end
				if(in == 412) begin
					state<=19;
					out<=78;
				end
				if(in == 413) begin
					state<=22;
					out<=79;
				end
				if(in == 414) begin
					state<=22;
					out<=80;
				end
				if(in == 415) begin
					state<=19;
					out<=81;
				end
				if(in == 416) begin
					state<=19;
					out<=82;
				end
				if(in == 417) begin
					state<=22;
					out<=83;
				end
				if(in == 418) begin
					state<=22;
					out<=84;
				end
				if(in == 419) begin
					state<=19;
					out<=85;
				end
				if(in == 420) begin
					state<=19;
					out<=86;
				end
				if(in == 421) begin
					state<=22;
					out<=87;
				end
				if(in == 422) begin
					state<=22;
					out<=88;
				end
				if(in == 423) begin
					state<=19;
					out<=89;
				end
				if(in == 424) begin
					state<=19;
					out<=90;
				end
				if(in == 425) begin
					state<=22;
					out<=91;
				end
				if(in == 426) begin
					state<=22;
					out<=92;
				end
				if(in == 427) begin
					state<=19;
					out<=93;
				end
				if(in == 428) begin
					state<=19;
					out<=94;
				end
				if(in == 429) begin
					state<=22;
					out<=95;
				end
				if(in == 430) begin
					state<=22;
					out<=96;
				end
				if(in == 431) begin
					state<=19;
					out<=97;
				end
				if(in == 432) begin
					state<=19;
					out<=98;
				end
				if(in == 433) begin
					state<=22;
					out<=99;
				end
				if(in == 434) begin
					state<=22;
					out<=100;
				end
				if(in == 435) begin
					state<=19;
					out<=101;
				end
				if(in == 436) begin
					state<=19;
					out<=102;
				end
				if(in == 437) begin
					state<=22;
					out<=103;
				end
				if(in == 438) begin
					state<=22;
					out<=104;
				end
				if(in == 439) begin
					state<=19;
					out<=105;
				end
				if(in == 440) begin
					state<=19;
					out<=106;
				end
				if(in == 441) begin
					state<=22;
					out<=107;
				end
				if(in == 442) begin
					state<=22;
					out<=108;
				end
				if(in == 443) begin
					state<=19;
					out<=109;
				end
				if(in == 444) begin
					state<=19;
					out<=110;
				end
				if(in == 445) begin
					state<=22;
					out<=111;
				end
				if(in == 446) begin
					state<=22;
					out<=112;
				end
				if(in == 447) begin
					state<=19;
					out<=113;
				end
				if(in == 448) begin
					state<=19;
					out<=114;
				end
				if(in == 449) begin
					state<=22;
					out<=115;
				end
				if(in == 450) begin
					state<=22;
					out<=116;
				end
				if(in == 451) begin
					state<=19;
					out<=117;
				end
				if(in == 452) begin
					state<=19;
					out<=118;
				end
				if(in == 453) begin
					state<=2;
					out<=119;
				end
				if(in == 454) begin
					state<=2;
					out<=120;
				end
				if(in == 455) begin
					state<=2;
					out<=121;
				end
				if(in == 456) begin
					state<=2;
					out<=122;
				end
				if(in == 457) begin
					state<=2;
					out<=123;
				end
				if(in == 458) begin
					state<=2;
					out<=124;
				end
				if(in == 459) begin
					state<=2;
					out<=125;
				end
				if(in == 460) begin
					state<=2;
					out<=126;
				end
				if(in == 461) begin
					state<=2;
					out<=127;
				end
				if(in == 462) begin
					state<=2;
					out<=128;
				end
				if(in == 463) begin
					state<=2;
					out<=129;
				end
				if(in == 464) begin
					state<=2;
					out<=130;
				end
				if(in == 465) begin
					state<=3;
					out<=131;
				end
				if(in == 466) begin
					state<=18;
					out<=132;
				end
				if(in == 467) begin
					state<=3;
					out<=133;
				end
				if(in == 468) begin
					state<=22;
					out<=134;
				end
				if(in == 469) begin
					state<=3;
					out<=135;
				end
				if(in == 470) begin
					state<=22;
					out<=136;
				end
				if(in == 471) begin
					state<=19;
					out<=137;
				end
				if(in == 472) begin
					state<=19;
					out<=138;
				end
				if(in == 473) begin
					state<=22;
					out<=139;
				end
				if(in == 474) begin
					state<=22;
					out<=140;
				end
				if(in == 475) begin
					state<=19;
					out<=141;
				end
				if(in == 476) begin
					state<=19;
					out<=142;
				end
				if(in == 477) begin
					state<=22;
					out<=143;
				end
				if(in == 478) begin
					state<=22;
					out<=144;
				end
				if(in == 479) begin
					state<=19;
					out<=145;
				end
				if(in == 480) begin
					state<=19;
					out<=146;
				end
				if(in == 481) begin
					state<=22;
					out<=147;
				end
				if(in == 482) begin
					state<=22;
					out<=148;
				end
				if(in == 483) begin
					state<=19;
					out<=149;
				end
				if(in == 484) begin
					state<=19;
					out<=150;
				end
				if(in == 485) begin
					state<=22;
					out<=151;
				end
				if(in == 486) begin
					state<=22;
					out<=152;
				end
				if(in == 487) begin
					state<=19;
					out<=153;
				end
				if(in == 488) begin
					state<=19;
					out<=154;
				end
				if(in == 489) begin
					state<=22;
					out<=155;
				end
				if(in == 490) begin
					state<=22;
					out<=156;
				end
				if(in == 491) begin
					state<=19;
					out<=157;
				end
				if(in == 492) begin
					state<=19;
					out<=158;
				end
				if(in == 493) begin
					state<=22;
					out<=159;
				end
				if(in == 494) begin
					state<=22;
					out<=160;
				end
				if(in == 495) begin
					state<=19;
					out<=161;
				end
				if(in == 496) begin
					state<=19;
					out<=162;
				end
				if(in == 497) begin
					state<=22;
					out<=163;
				end
				if(in == 498) begin
					state<=22;
					out<=164;
				end
				if(in == 499) begin
					state<=19;
					out<=165;
				end
				if(in == 500) begin
					state<=19;
					out<=166;
				end
				if(in == 501) begin
					state<=22;
					out<=167;
				end
				if(in == 502) begin
					state<=22;
					out<=168;
				end
				if(in == 503) begin
					state<=19;
					out<=169;
				end
				if(in == 504) begin
					state<=19;
					out<=170;
				end
				if(in == 505) begin
					state<=22;
					out<=171;
				end
				if(in == 506) begin
					state<=22;
					out<=172;
				end
				if(in == 507) begin
					state<=19;
					out<=173;
				end
				if(in == 508) begin
					state<=19;
					out<=174;
				end
				if(in == 509) begin
					state<=22;
					out<=175;
				end
				if(in == 510) begin
					state<=22;
					out<=176;
				end
				if(in == 511) begin
					state<=19;
					out<=177;
				end
				if(in == 512) begin
					state<=19;
					out<=178;
				end
				if(in == 513) begin
					state<=22;
					out<=179;
				end
				if(in == 514) begin
					state<=22;
					out<=180;
				end
				if(in == 515) begin
					state<=19;
					out<=181;
				end
				if(in == 516) begin
					state<=19;
					out<=182;
				end
				if(in == 517) begin
					state<=3;
					out<=183;
				end
				if(in == 518) begin
					state<=18;
					out<=184;
				end
				if(in == 519) begin
					state<=3;
					out<=185;
				end
				if(in == 520) begin
					state<=22;
					out<=186;
				end
				if(in == 521) begin
					state<=3;
					out<=187;
				end
				if(in == 522) begin
					state<=22;
					out<=188;
				end
				if(in == 523) begin
					state<=19;
					out<=189;
				end
				if(in == 524) begin
					state<=19;
					out<=190;
				end
				if(in == 525) begin
					state<=22;
					out<=191;
				end
				if(in == 526) begin
					state<=22;
					out<=192;
				end
				if(in == 527) begin
					state<=19;
					out<=193;
				end
				if(in == 528) begin
					state<=19;
					out<=194;
				end
				if(in == 529) begin
					state<=22;
					out<=195;
				end
				if(in == 530) begin
					state<=22;
					out<=196;
				end
				if(in == 531) begin
					state<=19;
					out<=197;
				end
				if(in == 532) begin
					state<=19;
					out<=198;
				end
				if(in == 533) begin
					state<=22;
					out<=199;
				end
				if(in == 534) begin
					state<=22;
					out<=200;
				end
				if(in == 535) begin
					state<=19;
					out<=201;
				end
				if(in == 536) begin
					state<=19;
					out<=202;
				end
				if(in == 537) begin
					state<=22;
					out<=203;
				end
				if(in == 538) begin
					state<=22;
					out<=204;
				end
				if(in == 539) begin
					state<=19;
					out<=205;
				end
				if(in == 540) begin
					state<=19;
					out<=206;
				end
				if(in == 541) begin
					state<=22;
					out<=207;
				end
				if(in == 542) begin
					state<=22;
					out<=208;
				end
				if(in == 543) begin
					state<=19;
					out<=209;
				end
				if(in == 544) begin
					state<=19;
					out<=210;
				end
				if(in == 545) begin
					state<=22;
					out<=211;
				end
				if(in == 546) begin
					state<=22;
					out<=212;
				end
				if(in == 547) begin
					state<=19;
					out<=213;
				end
				if(in == 548) begin
					state<=19;
					out<=214;
				end
				if(in == 549) begin
					state<=22;
					out<=215;
				end
				if(in == 550) begin
					state<=22;
					out<=216;
				end
				if(in == 551) begin
					state<=19;
					out<=217;
				end
				if(in == 552) begin
					state<=19;
					out<=218;
				end
				if(in == 553) begin
					state<=22;
					out<=219;
				end
				if(in == 554) begin
					state<=22;
					out<=220;
				end
				if(in == 555) begin
					state<=19;
					out<=221;
				end
				if(in == 556) begin
					state<=19;
					out<=222;
				end
				if(in == 557) begin
					state<=22;
					out<=223;
				end
				if(in == 558) begin
					state<=22;
					out<=224;
				end
				if(in == 559) begin
					state<=19;
					out<=225;
				end
				if(in == 560) begin
					state<=19;
					out<=226;
				end
				if(in == 561) begin
					state<=22;
					out<=227;
				end
				if(in == 562) begin
					state<=22;
					out<=228;
				end
				if(in == 563) begin
					state<=19;
					out<=229;
				end
				if(in == 564) begin
					state<=19;
					out<=230;
				end
				if(in == 565) begin
					state<=22;
					out<=231;
				end
				if(in == 566) begin
					state<=22;
					out<=232;
				end
				if(in == 567) begin
					state<=19;
					out<=233;
				end
				if(in == 568) begin
					state<=19;
					out<=234;
				end
				if(in == 569) begin
					state<=2;
					out<=235;
				end
				if(in == 570) begin
					state<=2;
					out<=236;
				end
				if(in == 571) begin
					state<=2;
					out<=237;
				end
				if(in == 572) begin
					state<=2;
					out<=238;
				end
				if(in == 573) begin
					state<=2;
					out<=239;
				end
				if(in == 574) begin
					state<=2;
					out<=240;
				end
				if(in == 575) begin
					state<=2;
					out<=241;
				end
				if(in == 576) begin
					state<=2;
					out<=242;
				end
				if(in == 577) begin
					state<=2;
					out<=243;
				end
				if(in == 578) begin
					state<=2;
					out<=244;
				end
				if(in == 579) begin
					state<=2;
					out<=245;
				end
				if(in == 580) begin
					state<=2;
					out<=246;
				end
				if(in == 581) begin
					state<=3;
					out<=247;
				end
				if(in == 582) begin
					state<=18;
					out<=248;
				end
				if(in == 583) begin
					state<=3;
					out<=249;
				end
				if(in == 584) begin
					state<=22;
					out<=250;
				end
				if(in == 585) begin
					state<=3;
					out<=251;
				end
				if(in == 586) begin
					state<=22;
					out<=252;
				end
				if(in == 587) begin
					state<=19;
					out<=253;
				end
				if(in == 588) begin
					state<=19;
					out<=254;
				end
				if(in == 589) begin
					state<=22;
					out<=255;
				end
				if(in == 590) begin
					state<=22;
					out<=0;
				end
				if(in == 591) begin
					state<=19;
					out<=1;
				end
				if(in == 592) begin
					state<=19;
					out<=2;
				end
				if(in == 593) begin
					state<=22;
					out<=3;
				end
				if(in == 594) begin
					state<=22;
					out<=4;
				end
				if(in == 595) begin
					state<=19;
					out<=5;
				end
				if(in == 596) begin
					state<=19;
					out<=6;
				end
				if(in == 597) begin
					state<=22;
					out<=7;
				end
				if(in == 598) begin
					state<=22;
					out<=8;
				end
				if(in == 599) begin
					state<=19;
					out<=9;
				end
				if(in == 600) begin
					state<=19;
					out<=10;
				end
				if(in == 601) begin
					state<=22;
					out<=11;
				end
				if(in == 602) begin
					state<=22;
					out<=12;
				end
				if(in == 603) begin
					state<=19;
					out<=13;
				end
				if(in == 604) begin
					state<=19;
					out<=14;
				end
				if(in == 605) begin
					state<=22;
					out<=15;
				end
				if(in == 606) begin
					state<=22;
					out<=16;
				end
				if(in == 607) begin
					state<=19;
					out<=17;
				end
				if(in == 608) begin
					state<=19;
					out<=18;
				end
				if(in == 609) begin
					state<=22;
					out<=19;
				end
				if(in == 610) begin
					state<=22;
					out<=20;
				end
				if(in == 611) begin
					state<=19;
					out<=21;
				end
				if(in == 612) begin
					state<=19;
					out<=22;
				end
				if(in == 613) begin
					state<=22;
					out<=23;
				end
				if(in == 614) begin
					state<=22;
					out<=24;
				end
				if(in == 615) begin
					state<=19;
					out<=25;
				end
				if(in == 616) begin
					state<=19;
					out<=26;
				end
				if(in == 617) begin
					state<=22;
					out<=27;
				end
				if(in == 618) begin
					state<=22;
					out<=28;
				end
				if(in == 619) begin
					state<=19;
					out<=29;
				end
				if(in == 620) begin
					state<=19;
					out<=30;
				end
				if(in == 621) begin
					state<=22;
					out<=31;
				end
				if(in == 622) begin
					state<=22;
					out<=32;
				end
				if(in == 623) begin
					state<=19;
					out<=33;
				end
				if(in == 624) begin
					state<=19;
					out<=34;
				end
				if(in == 625) begin
					state<=22;
					out<=35;
				end
				if(in == 626) begin
					state<=22;
					out<=36;
				end
				if(in == 627) begin
					state<=19;
					out<=37;
				end
				if(in == 628) begin
					state<=19;
					out<=38;
				end
				if(in == 629) begin
					state<=22;
					out<=39;
				end
				if(in == 630) begin
					state<=22;
					out<=40;
				end
				if(in == 631) begin
					state<=19;
					out<=41;
				end
				if(in == 632) begin
					state<=19;
					out<=42;
				end
				if(in == 633) begin
					state<=3;
					out<=43;
				end
				if(in == 634) begin
					state<=18;
					out<=44;
				end
				if(in == 635) begin
					state<=3;
					out<=45;
				end
				if(in == 636) begin
					state<=22;
					out<=46;
				end
				if(in == 637) begin
					state<=3;
					out<=47;
				end
				if(in == 638) begin
					state<=22;
					out<=48;
				end
				if(in == 639) begin
					state<=19;
					out<=49;
				end
				if(in == 640) begin
					state<=19;
					out<=50;
				end
				if(in == 641) begin
					state<=22;
					out<=51;
				end
				if(in == 642) begin
					state<=22;
					out<=52;
				end
				if(in == 643) begin
					state<=19;
					out<=53;
				end
				if(in == 644) begin
					state<=19;
					out<=54;
				end
				if(in == 645) begin
					state<=22;
					out<=55;
				end
				if(in == 646) begin
					state<=22;
					out<=56;
				end
				if(in == 647) begin
					state<=19;
					out<=57;
				end
				if(in == 648) begin
					state<=19;
					out<=58;
				end
				if(in == 649) begin
					state<=22;
					out<=59;
				end
				if(in == 650) begin
					state<=22;
					out<=60;
				end
				if(in == 651) begin
					state<=19;
					out<=61;
				end
				if(in == 652) begin
					state<=19;
					out<=62;
				end
				if(in == 653) begin
					state<=22;
					out<=63;
				end
				if(in == 654) begin
					state<=22;
					out<=64;
				end
				if(in == 655) begin
					state<=19;
					out<=65;
				end
				if(in == 656) begin
					state<=19;
					out<=66;
				end
				if(in == 657) begin
					state<=22;
					out<=67;
				end
				if(in == 658) begin
					state<=22;
					out<=68;
				end
				if(in == 659) begin
					state<=19;
					out<=69;
				end
				if(in == 660) begin
					state<=19;
					out<=70;
				end
				if(in == 661) begin
					state<=22;
					out<=71;
				end
				if(in == 662) begin
					state<=22;
					out<=72;
				end
				if(in == 663) begin
					state<=19;
					out<=73;
				end
				if(in == 664) begin
					state<=19;
					out<=74;
				end
				if(in == 665) begin
					state<=22;
					out<=75;
				end
				if(in == 666) begin
					state<=22;
					out<=76;
				end
				if(in == 667) begin
					state<=19;
					out<=77;
				end
				if(in == 668) begin
					state<=19;
					out<=78;
				end
				if(in == 669) begin
					state<=22;
					out<=79;
				end
				if(in == 670) begin
					state<=22;
					out<=80;
				end
				if(in == 671) begin
					state<=19;
					out<=81;
				end
				if(in == 672) begin
					state<=19;
					out<=82;
				end
				if(in == 673) begin
					state<=22;
					out<=83;
				end
				if(in == 674) begin
					state<=22;
					out<=84;
				end
				if(in == 675) begin
					state<=19;
					out<=85;
				end
				if(in == 676) begin
					state<=19;
					out<=86;
				end
				if(in == 677) begin
					state<=22;
					out<=87;
				end
				if(in == 678) begin
					state<=22;
					out<=88;
				end
				if(in == 679) begin
					state<=19;
					out<=89;
				end
				if(in == 680) begin
					state<=19;
					out<=90;
				end
				if(in == 681) begin
					state<=22;
					out<=91;
				end
				if(in == 682) begin
					state<=22;
					out<=92;
				end
				if(in == 683) begin
					state<=19;
					out<=93;
				end
				if(in == 684) begin
					state<=19;
					out<=94;
				end
				if(in == 685) begin
					state<=2;
					out<=95;
				end
				if(in == 686) begin
					state<=2;
					out<=96;
				end
				if(in == 687) begin
					state<=2;
					out<=97;
				end
				if(in == 688) begin
					state<=2;
					out<=98;
				end
				if(in == 689) begin
					state<=2;
					out<=99;
				end
				if(in == 690) begin
					state<=2;
					out<=100;
				end
				if(in == 691) begin
					state<=2;
					out<=101;
				end
				if(in == 692) begin
					state<=2;
					out<=102;
				end
				if(in == 693) begin
					state<=2;
					out<=103;
				end
				if(in == 694) begin
					state<=2;
					out<=104;
				end
				if(in == 695) begin
					state<=2;
					out<=105;
				end
				if(in == 696) begin
					state<=2;
					out<=106;
				end
				if(in == 697) begin
					state<=3;
					out<=107;
				end
				if(in == 698) begin
					state<=18;
					out<=108;
				end
				if(in == 699) begin
					state<=3;
					out<=109;
				end
				if(in == 700) begin
					state<=22;
					out<=110;
				end
				if(in == 701) begin
					state<=3;
					out<=111;
				end
				if(in == 702) begin
					state<=22;
					out<=112;
				end
				if(in == 703) begin
					state<=19;
					out<=113;
				end
				if(in == 704) begin
					state<=19;
					out<=114;
				end
				if(in == 705) begin
					state<=22;
					out<=115;
				end
				if(in == 706) begin
					state<=22;
					out<=116;
				end
				if(in == 707) begin
					state<=19;
					out<=117;
				end
				if(in == 708) begin
					state<=19;
					out<=118;
				end
				if(in == 709) begin
					state<=22;
					out<=119;
				end
				if(in == 710) begin
					state<=22;
					out<=120;
				end
				if(in == 711) begin
					state<=19;
					out<=121;
				end
				if(in == 712) begin
					state<=19;
					out<=122;
				end
				if(in == 713) begin
					state<=22;
					out<=123;
				end
				if(in == 714) begin
					state<=22;
					out<=124;
				end
				if(in == 715) begin
					state<=19;
					out<=125;
				end
				if(in == 716) begin
					state<=19;
					out<=126;
				end
				if(in == 717) begin
					state<=22;
					out<=127;
				end
				if(in == 718) begin
					state<=22;
					out<=128;
				end
				if(in == 719) begin
					state<=19;
					out<=129;
				end
				if(in == 720) begin
					state<=19;
					out<=130;
				end
				if(in == 721) begin
					state<=22;
					out<=131;
				end
				if(in == 722) begin
					state<=22;
					out<=132;
				end
				if(in == 723) begin
					state<=19;
					out<=133;
				end
				if(in == 724) begin
					state<=19;
					out<=134;
				end
				if(in == 725) begin
					state<=22;
					out<=135;
				end
				if(in == 726) begin
					state<=22;
					out<=136;
				end
				if(in == 727) begin
					state<=19;
					out<=137;
				end
				if(in == 728) begin
					state<=19;
					out<=138;
				end
				if(in == 729) begin
					state<=22;
					out<=139;
				end
				if(in == 730) begin
					state<=22;
					out<=140;
				end
				if(in == 731) begin
					state<=19;
					out<=141;
				end
				if(in == 732) begin
					state<=19;
					out<=142;
				end
				if(in == 733) begin
					state<=22;
					out<=143;
				end
				if(in == 734) begin
					state<=22;
					out<=144;
				end
				if(in == 735) begin
					state<=19;
					out<=145;
				end
				if(in == 736) begin
					state<=19;
					out<=146;
				end
				if(in == 737) begin
					state<=22;
					out<=147;
				end
				if(in == 738) begin
					state<=22;
					out<=148;
				end
				if(in == 739) begin
					state<=19;
					out<=149;
				end
				if(in == 740) begin
					state<=19;
					out<=150;
				end
				if(in == 741) begin
					state<=22;
					out<=151;
				end
				if(in == 742) begin
					state<=22;
					out<=152;
				end
				if(in == 743) begin
					state<=19;
					out<=153;
				end
				if(in == 744) begin
					state<=19;
					out<=154;
				end
				if(in == 745) begin
					state<=22;
					out<=155;
				end
				if(in == 746) begin
					state<=22;
					out<=156;
				end
				if(in == 747) begin
					state<=19;
					out<=157;
				end
				if(in == 748) begin
					state<=19;
					out<=158;
				end
				if(in == 749) begin
					state<=3;
					out<=159;
				end
				if(in == 750) begin
					state<=18;
					out<=160;
				end
				if(in == 751) begin
					state<=3;
					out<=161;
				end
				if(in == 752) begin
					state<=22;
					out<=162;
				end
				if(in == 753) begin
					state<=3;
					out<=163;
				end
				if(in == 754) begin
					state<=22;
					out<=164;
				end
				if(in == 755) begin
					state<=19;
					out<=165;
				end
				if(in == 756) begin
					state<=19;
					out<=166;
				end
				if(in == 757) begin
					state<=22;
					out<=167;
				end
				if(in == 758) begin
					state<=22;
					out<=168;
				end
				if(in == 759) begin
					state<=19;
					out<=169;
				end
				if(in == 760) begin
					state<=19;
					out<=170;
				end
				if(in == 761) begin
					state<=22;
					out<=171;
				end
				if(in == 762) begin
					state<=22;
					out<=172;
				end
				if(in == 763) begin
					state<=19;
					out<=173;
				end
				if(in == 764) begin
					state<=19;
					out<=174;
				end
				if(in == 765) begin
					state<=22;
					out<=175;
				end
				if(in == 766) begin
					state<=22;
					out<=176;
				end
				if(in == 767) begin
					state<=19;
					out<=177;
				end
				if(in == 768) begin
					state<=19;
					out<=178;
				end
				if(in == 769) begin
					state<=22;
					out<=179;
				end
				if(in == 770) begin
					state<=22;
					out<=180;
				end
				if(in == 771) begin
					state<=19;
					out<=181;
				end
				if(in == 772) begin
					state<=19;
					out<=182;
				end
				if(in == 773) begin
					state<=22;
					out<=183;
				end
				if(in == 774) begin
					state<=22;
					out<=184;
				end
				if(in == 775) begin
					state<=19;
					out<=185;
				end
				if(in == 776) begin
					state<=19;
					out<=186;
				end
				if(in == 777) begin
					state<=22;
					out<=187;
				end
				if(in == 778) begin
					state<=22;
					out<=188;
				end
				if(in == 779) begin
					state<=19;
					out<=189;
				end
				if(in == 780) begin
					state<=19;
					out<=190;
				end
				if(in == 781) begin
					state<=22;
					out<=191;
				end
				if(in == 782) begin
					state<=22;
					out<=192;
				end
				if(in == 783) begin
					state<=19;
					out<=193;
				end
				if(in == 784) begin
					state<=19;
					out<=194;
				end
				if(in == 785) begin
					state<=22;
					out<=195;
				end
				if(in == 786) begin
					state<=22;
					out<=196;
				end
				if(in == 787) begin
					state<=19;
					out<=197;
				end
				if(in == 788) begin
					state<=19;
					out<=198;
				end
				if(in == 789) begin
					state<=22;
					out<=199;
				end
				if(in == 790) begin
					state<=22;
					out<=200;
				end
				if(in == 791) begin
					state<=19;
					out<=201;
				end
				if(in == 792) begin
					state<=19;
					out<=202;
				end
				if(in == 793) begin
					state<=22;
					out<=203;
				end
				if(in == 794) begin
					state<=22;
					out<=204;
				end
				if(in == 795) begin
					state<=19;
					out<=205;
				end
				if(in == 796) begin
					state<=19;
					out<=206;
				end
				if(in == 797) begin
					state<=22;
					out<=207;
				end
				if(in == 798) begin
					state<=22;
					out<=208;
				end
				if(in == 799) begin
					state<=19;
					out<=209;
				end
				if(in == 800) begin
					state<=19;
					out<=210;
				end
				if(in == 801) begin
					state<=2;
					out<=211;
				end
				if(in == 802) begin
					state<=2;
					out<=212;
				end
				if(in == 803) begin
					state<=2;
					out<=213;
				end
				if(in == 804) begin
					state<=2;
					out<=214;
				end
				if(in == 805) begin
					state<=2;
					out<=215;
				end
				if(in == 806) begin
					state<=2;
					out<=216;
				end
				if(in == 807) begin
					state<=2;
					out<=217;
				end
				if(in == 808) begin
					state<=2;
					out<=218;
				end
				if(in == 809) begin
					state<=2;
					out<=219;
				end
				if(in == 810) begin
					state<=2;
					out<=220;
				end
				if(in == 811) begin
					state<=2;
					out<=221;
				end
				if(in == 812) begin
					state<=2;
					out<=222;
				end
				if(in == 813) begin
					state<=3;
					out<=223;
				end
				if(in == 814) begin
					state<=18;
					out<=224;
				end
				if(in == 815) begin
					state<=3;
					out<=225;
				end
				if(in == 816) begin
					state<=22;
					out<=226;
				end
				if(in == 817) begin
					state<=3;
					out<=227;
				end
				if(in == 818) begin
					state<=22;
					out<=228;
				end
				if(in == 819) begin
					state<=19;
					out<=229;
				end
				if(in == 820) begin
					state<=19;
					out<=230;
				end
				if(in == 821) begin
					state<=22;
					out<=231;
				end
				if(in == 822) begin
					state<=22;
					out<=232;
				end
				if(in == 823) begin
					state<=19;
					out<=233;
				end
				if(in == 824) begin
					state<=19;
					out<=234;
				end
				if(in == 825) begin
					state<=22;
					out<=235;
				end
				if(in == 826) begin
					state<=22;
					out<=236;
				end
				if(in == 827) begin
					state<=19;
					out<=237;
				end
				if(in == 828) begin
					state<=19;
					out<=238;
				end
				if(in == 829) begin
					state<=22;
					out<=239;
				end
				if(in == 830) begin
					state<=22;
					out<=240;
				end
				if(in == 831) begin
					state<=19;
					out<=241;
				end
				if(in == 832) begin
					state<=19;
					out<=242;
				end
				if(in == 833) begin
					state<=22;
					out<=243;
				end
				if(in == 834) begin
					state<=22;
					out<=244;
				end
				if(in == 835) begin
					state<=19;
					out<=245;
				end
				if(in == 836) begin
					state<=19;
					out<=246;
				end
				if(in == 837) begin
					state<=22;
					out<=247;
				end
				if(in == 838) begin
					state<=22;
					out<=248;
				end
				if(in == 839) begin
					state<=19;
					out<=249;
				end
				if(in == 840) begin
					state<=19;
					out<=250;
				end
				if(in == 841) begin
					state<=22;
					out<=251;
				end
				if(in == 842) begin
					state<=22;
					out<=252;
				end
				if(in == 843) begin
					state<=19;
					out<=253;
				end
				if(in == 844) begin
					state<=19;
					out<=254;
				end
				if(in == 845) begin
					state<=22;
					out<=255;
				end
				if(in == 846) begin
					state<=22;
					out<=0;
				end
				if(in == 847) begin
					state<=19;
					out<=1;
				end
				if(in == 848) begin
					state<=19;
					out<=2;
				end
				if(in == 849) begin
					state<=22;
					out<=3;
				end
				if(in == 850) begin
					state<=22;
					out<=4;
				end
				if(in == 851) begin
					state<=19;
					out<=5;
				end
				if(in == 852) begin
					state<=19;
					out<=6;
				end
				if(in == 853) begin
					state<=22;
					out<=7;
				end
				if(in == 854) begin
					state<=22;
					out<=8;
				end
				if(in == 855) begin
					state<=19;
					out<=9;
				end
				if(in == 856) begin
					state<=19;
					out<=10;
				end
				if(in == 857) begin
					state<=22;
					out<=11;
				end
				if(in == 858) begin
					state<=22;
					out<=12;
				end
				if(in == 859) begin
					state<=19;
					out<=13;
				end
				if(in == 860) begin
					state<=19;
					out<=14;
				end
				if(in == 861) begin
					state<=22;
					out<=15;
				end
				if(in == 862) begin
					state<=22;
					out<=16;
				end
				if(in == 863) begin
					state<=19;
					out<=17;
				end
				if(in == 864) begin
					state<=19;
					out<=18;
				end
				if(in == 865) begin
					state<=3;
					out<=19;
				end
				if(in == 866) begin
					state<=18;
					out<=20;
				end
				if(in == 867) begin
					state<=3;
					out<=21;
				end
				if(in == 868) begin
					state<=22;
					out<=22;
				end
				if(in == 869) begin
					state<=3;
					out<=23;
				end
				if(in == 870) begin
					state<=22;
					out<=24;
				end
				if(in == 871) begin
					state<=19;
					out<=25;
				end
				if(in == 872) begin
					state<=19;
					out<=26;
				end
				if(in == 873) begin
					state<=22;
					out<=27;
				end
				if(in == 874) begin
					state<=22;
					out<=28;
				end
				if(in == 875) begin
					state<=19;
					out<=29;
				end
				if(in == 876) begin
					state<=19;
					out<=30;
				end
				if(in == 877) begin
					state<=22;
					out<=31;
				end
				if(in == 878) begin
					state<=22;
					out<=32;
				end
				if(in == 879) begin
					state<=19;
					out<=33;
				end
				if(in == 880) begin
					state<=19;
					out<=34;
				end
				if(in == 881) begin
					state<=22;
					out<=35;
				end
				if(in == 882) begin
					state<=22;
					out<=36;
				end
				if(in == 883) begin
					state<=19;
					out<=37;
				end
				if(in == 884) begin
					state<=19;
					out<=38;
				end
				if(in == 885) begin
					state<=22;
					out<=39;
				end
				if(in == 886) begin
					state<=22;
					out<=40;
				end
				if(in == 887) begin
					state<=19;
					out<=41;
				end
				if(in == 888) begin
					state<=19;
					out<=42;
				end
				if(in == 889) begin
					state<=22;
					out<=43;
				end
				if(in == 890) begin
					state<=22;
					out<=44;
				end
				if(in == 891) begin
					state<=19;
					out<=45;
				end
				if(in == 892) begin
					state<=19;
					out<=46;
				end
				if(in == 893) begin
					state<=22;
					out<=47;
				end
				if(in == 894) begin
					state<=22;
					out<=48;
				end
				if(in == 895) begin
					state<=19;
					out<=49;
				end
				if(in == 896) begin
					state<=19;
					out<=50;
				end
				if(in == 897) begin
					state<=22;
					out<=51;
				end
				if(in == 898) begin
					state<=22;
					out<=52;
				end
				if(in == 899) begin
					state<=19;
					out<=53;
				end
				if(in == 900) begin
					state<=19;
					out<=54;
				end
				if(in == 901) begin
					state<=22;
					out<=55;
				end
				if(in == 902) begin
					state<=22;
					out<=56;
				end
				if(in == 903) begin
					state<=19;
					out<=57;
				end
				if(in == 904) begin
					state<=19;
					out<=58;
				end
				if(in == 905) begin
					state<=22;
					out<=59;
				end
				if(in == 906) begin
					state<=22;
					out<=60;
				end
				if(in == 907) begin
					state<=19;
					out<=61;
				end
				if(in == 908) begin
					state<=19;
					out<=62;
				end
				if(in == 909) begin
					state<=22;
					out<=63;
				end
				if(in == 910) begin
					state<=22;
					out<=64;
				end
				if(in == 911) begin
					state<=19;
					out<=65;
				end
				if(in == 912) begin
					state<=19;
					out<=66;
				end
				if(in == 913) begin
					state<=22;
					out<=67;
				end
				if(in == 914) begin
					state<=22;
					out<=68;
				end
				if(in == 915) begin
					state<=19;
					out<=69;
				end
				if(in == 916) begin
					state<=19;
					out<=70;
				end
				if(in == 917) begin
					state<=2;
					out<=71;
				end
				if(in == 918) begin
					state<=2;
					out<=72;
				end
				if(in == 919) begin
					state<=2;
					out<=73;
				end
				if(in == 920) begin
					state<=2;
					out<=74;
				end
				if(in == 921) begin
					state<=2;
					out<=75;
				end
				if(in == 922) begin
					state<=2;
					out<=76;
				end
				if(in == 923) begin
					state<=2;
					out<=77;
				end
				if(in == 924) begin
					state<=2;
					out<=78;
				end
				if(in == 925) begin
					state<=2;
					out<=79;
				end
				if(in == 926) begin
					state<=2;
					out<=80;
				end
				if(in == 927) begin
					state<=2;
					out<=81;
				end
				if(in == 928) begin
					state<=2;
					out<=82;
				end
			end
			19: begin
				if(in == 0) begin
					state<=3;
					out<=83;
				end
				if(in == 1) begin
					state<=1;
					out<=84;
				end
				if(in == 2) begin
					state<=19;
					out<=85;
				end
				if(in == 3) begin
					state<=3;
					out<=86;
				end
				if(in == 4) begin
					state<=20;
					out<=87;
				end
				if(in == 5) begin
					state<=3;
					out<=88;
				end
				if(in == 6) begin
					state<=20;
					out<=89;
				end
				if(in == 7) begin
					state<=20;
					out<=90;
				end
				if(in == 8) begin
					state<=20;
					out<=91;
				end
				if(in == 9) begin
					state<=20;
					out<=92;
				end
				if(in == 10) begin
					state<=20;
					out<=93;
				end
				if(in == 11) begin
					state<=20;
					out<=94;
				end
				if(in == 12) begin
					state<=20;
					out<=95;
				end
				if(in == 13) begin
					state<=20;
					out<=96;
				end
				if(in == 14) begin
					state<=20;
					out<=97;
				end
				if(in == 15) begin
					state<=20;
					out<=98;
				end
				if(in == 16) begin
					state<=20;
					out<=99;
				end
				if(in == 17) begin
					state<=20;
					out<=100;
				end
				if(in == 18) begin
					state<=20;
					out<=101;
				end
				if(in == 19) begin
					state<=20;
					out<=102;
				end
				if(in == 20) begin
					state<=20;
					out<=103;
				end
				if(in == 21) begin
					state<=20;
					out<=104;
				end
				if(in == 22) begin
					state<=20;
					out<=105;
				end
				if(in == 23) begin
					state<=20;
					out<=106;
				end
				if(in == 24) begin
					state<=20;
					out<=107;
				end
				if(in == 25) begin
					state<=20;
					out<=108;
				end
				if(in == 26) begin
					state<=20;
					out<=109;
				end
				if(in == 27) begin
					state<=20;
					out<=110;
				end
				if(in == 28) begin
					state<=20;
					out<=111;
				end
				if(in == 29) begin
					state<=20;
					out<=112;
				end
				if(in == 30) begin
					state<=20;
					out<=113;
				end
				if(in == 31) begin
					state<=20;
					out<=114;
				end
				if(in == 32) begin
					state<=20;
					out<=115;
				end
				if(in == 33) begin
					state<=20;
					out<=116;
				end
				if(in == 34) begin
					state<=20;
					out<=117;
				end
				if(in == 35) begin
					state<=20;
					out<=118;
				end
				if(in == 36) begin
					state<=20;
					out<=119;
				end
				if(in == 37) begin
					state<=20;
					out<=120;
				end
				if(in == 38) begin
					state<=20;
					out<=121;
				end
				if(in == 39) begin
					state<=20;
					out<=122;
				end
				if(in == 40) begin
					state<=20;
					out<=123;
				end
				if(in == 41) begin
					state<=20;
					out<=124;
				end
				if(in == 42) begin
					state<=20;
					out<=125;
				end
				if(in == 43) begin
					state<=20;
					out<=126;
				end
				if(in == 44) begin
					state<=20;
					out<=127;
				end
				if(in == 45) begin
					state<=20;
					out<=128;
				end
				if(in == 46) begin
					state<=20;
					out<=129;
				end
				if(in == 47) begin
					state<=20;
					out<=130;
				end
				if(in == 48) begin
					state<=20;
					out<=131;
				end
				if(in == 49) begin
					state<=20;
					out<=132;
				end
				if(in == 50) begin
					state<=20;
					out<=133;
				end
				if(in == 51) begin
					state<=20;
					out<=134;
				end
				if(in == 52) begin
					state<=20;
					out<=135;
				end
				if(in == 53) begin
					state<=3;
					out<=136;
				end
				if(in == 54) begin
					state<=19;
					out<=137;
				end
				if(in == 55) begin
					state<=3;
					out<=138;
				end
				if(in == 56) begin
					state<=20;
					out<=139;
				end
				if(in == 57) begin
					state<=3;
					out<=140;
				end
				if(in == 58) begin
					state<=20;
					out<=141;
				end
				if(in == 59) begin
					state<=20;
					out<=142;
				end
				if(in == 60) begin
					state<=20;
					out<=143;
				end
				if(in == 61) begin
					state<=20;
					out<=144;
				end
				if(in == 62) begin
					state<=20;
					out<=145;
				end
				if(in == 63) begin
					state<=20;
					out<=146;
				end
				if(in == 64) begin
					state<=20;
					out<=147;
				end
				if(in == 65) begin
					state<=20;
					out<=148;
				end
				if(in == 66) begin
					state<=20;
					out<=149;
				end
				if(in == 67) begin
					state<=20;
					out<=150;
				end
				if(in == 68) begin
					state<=20;
					out<=151;
				end
				if(in == 69) begin
					state<=20;
					out<=152;
				end
				if(in == 70) begin
					state<=20;
					out<=153;
				end
				if(in == 71) begin
					state<=20;
					out<=154;
				end
				if(in == 72) begin
					state<=20;
					out<=155;
				end
				if(in == 73) begin
					state<=20;
					out<=156;
				end
				if(in == 74) begin
					state<=20;
					out<=157;
				end
				if(in == 75) begin
					state<=20;
					out<=158;
				end
				if(in == 76) begin
					state<=20;
					out<=159;
				end
				if(in == 77) begin
					state<=20;
					out<=160;
				end
				if(in == 78) begin
					state<=20;
					out<=161;
				end
				if(in == 79) begin
					state<=20;
					out<=162;
				end
				if(in == 80) begin
					state<=20;
					out<=163;
				end
				if(in == 81) begin
					state<=20;
					out<=164;
				end
				if(in == 82) begin
					state<=20;
					out<=165;
				end
				if(in == 83) begin
					state<=20;
					out<=166;
				end
				if(in == 84) begin
					state<=20;
					out<=167;
				end
				if(in == 85) begin
					state<=20;
					out<=168;
				end
				if(in == 86) begin
					state<=20;
					out<=169;
				end
				if(in == 87) begin
					state<=20;
					out<=170;
				end
				if(in == 88) begin
					state<=20;
					out<=171;
				end
				if(in == 89) begin
					state<=20;
					out<=172;
				end
				if(in == 90) begin
					state<=20;
					out<=173;
				end
				if(in == 91) begin
					state<=20;
					out<=174;
				end
				if(in == 92) begin
					state<=20;
					out<=175;
				end
				if(in == 93) begin
					state<=20;
					out<=176;
				end
				if(in == 94) begin
					state<=20;
					out<=177;
				end
				if(in == 95) begin
					state<=20;
					out<=178;
				end
				if(in == 96) begin
					state<=20;
					out<=179;
				end
				if(in == 97) begin
					state<=20;
					out<=180;
				end
				if(in == 98) begin
					state<=20;
					out<=181;
				end
				if(in == 99) begin
					state<=20;
					out<=182;
				end
				if(in == 100) begin
					state<=20;
					out<=183;
				end
				if(in == 101) begin
					state<=20;
					out<=184;
				end
				if(in == 102) begin
					state<=20;
					out<=185;
				end
				if(in == 103) begin
					state<=20;
					out<=186;
				end
				if(in == 104) begin
					state<=20;
					out<=187;
				end
				if(in == 105) begin
					state<=2;
					out<=188;
				end
				if(in == 106) begin
					state<=2;
					out<=189;
				end
				if(in == 107) begin
					state<=2;
					out<=190;
				end
				if(in == 108) begin
					state<=2;
					out<=191;
				end
				if(in == 109) begin
					state<=2;
					out<=192;
				end
				if(in == 110) begin
					state<=2;
					out<=193;
				end
				if(in == 111) begin
					state<=2;
					out<=194;
				end
				if(in == 112) begin
					state<=2;
					out<=195;
				end
				if(in == 113) begin
					state<=2;
					out<=196;
				end
				if(in == 114) begin
					state<=2;
					out<=197;
				end
				if(in == 115) begin
					state<=2;
					out<=198;
				end
				if(in == 116) begin
					state<=2;
					out<=199;
				end
				if(in == 117) begin
					state<=3;
					out<=200;
				end
				if(in == 118) begin
					state<=19;
					out<=201;
				end
				if(in == 119) begin
					state<=3;
					out<=202;
				end
				if(in == 120) begin
					state<=20;
					out<=203;
				end
				if(in == 121) begin
					state<=3;
					out<=204;
				end
				if(in == 122) begin
					state<=20;
					out<=205;
				end
				if(in == 123) begin
					state<=20;
					out<=206;
				end
				if(in == 124) begin
					state<=20;
					out<=207;
				end
				if(in == 125) begin
					state<=20;
					out<=208;
				end
				if(in == 126) begin
					state<=20;
					out<=209;
				end
				if(in == 127) begin
					state<=20;
					out<=210;
				end
				if(in == 128) begin
					state<=20;
					out<=211;
				end
				if(in == 129) begin
					state<=20;
					out<=212;
				end
				if(in == 130) begin
					state<=20;
					out<=213;
				end
				if(in == 131) begin
					state<=20;
					out<=214;
				end
				if(in == 132) begin
					state<=20;
					out<=215;
				end
				if(in == 133) begin
					state<=20;
					out<=216;
				end
				if(in == 134) begin
					state<=20;
					out<=217;
				end
				if(in == 135) begin
					state<=20;
					out<=218;
				end
				if(in == 136) begin
					state<=20;
					out<=219;
				end
				if(in == 137) begin
					state<=20;
					out<=220;
				end
				if(in == 138) begin
					state<=20;
					out<=221;
				end
				if(in == 139) begin
					state<=20;
					out<=222;
				end
				if(in == 140) begin
					state<=20;
					out<=223;
				end
				if(in == 141) begin
					state<=20;
					out<=224;
				end
				if(in == 142) begin
					state<=20;
					out<=225;
				end
				if(in == 143) begin
					state<=20;
					out<=226;
				end
				if(in == 144) begin
					state<=20;
					out<=227;
				end
				if(in == 145) begin
					state<=20;
					out<=228;
				end
				if(in == 146) begin
					state<=20;
					out<=229;
				end
				if(in == 147) begin
					state<=20;
					out<=230;
				end
				if(in == 148) begin
					state<=20;
					out<=231;
				end
				if(in == 149) begin
					state<=20;
					out<=232;
				end
				if(in == 150) begin
					state<=20;
					out<=233;
				end
				if(in == 151) begin
					state<=20;
					out<=234;
				end
				if(in == 152) begin
					state<=20;
					out<=235;
				end
				if(in == 153) begin
					state<=20;
					out<=236;
				end
				if(in == 154) begin
					state<=20;
					out<=237;
				end
				if(in == 155) begin
					state<=20;
					out<=238;
				end
				if(in == 156) begin
					state<=20;
					out<=239;
				end
				if(in == 157) begin
					state<=20;
					out<=240;
				end
				if(in == 158) begin
					state<=20;
					out<=241;
				end
				if(in == 159) begin
					state<=20;
					out<=242;
				end
				if(in == 160) begin
					state<=20;
					out<=243;
				end
				if(in == 161) begin
					state<=20;
					out<=244;
				end
				if(in == 162) begin
					state<=20;
					out<=245;
				end
				if(in == 163) begin
					state<=20;
					out<=246;
				end
				if(in == 164) begin
					state<=20;
					out<=247;
				end
				if(in == 165) begin
					state<=20;
					out<=248;
				end
				if(in == 166) begin
					state<=20;
					out<=249;
				end
				if(in == 167) begin
					state<=20;
					out<=250;
				end
				if(in == 168) begin
					state<=20;
					out<=251;
				end
				if(in == 169) begin
					state<=3;
					out<=252;
				end
				if(in == 170) begin
					state<=19;
					out<=253;
				end
				if(in == 171) begin
					state<=3;
					out<=254;
				end
				if(in == 172) begin
					state<=20;
					out<=255;
				end
				if(in == 173) begin
					state<=3;
					out<=0;
				end
				if(in == 174) begin
					state<=20;
					out<=1;
				end
				if(in == 175) begin
					state<=20;
					out<=2;
				end
				if(in == 176) begin
					state<=20;
					out<=3;
				end
				if(in == 177) begin
					state<=20;
					out<=4;
				end
				if(in == 178) begin
					state<=20;
					out<=5;
				end
				if(in == 179) begin
					state<=20;
					out<=6;
				end
				if(in == 180) begin
					state<=20;
					out<=7;
				end
				if(in == 181) begin
					state<=20;
					out<=8;
				end
				if(in == 182) begin
					state<=20;
					out<=9;
				end
				if(in == 183) begin
					state<=20;
					out<=10;
				end
				if(in == 184) begin
					state<=20;
					out<=11;
				end
				if(in == 185) begin
					state<=20;
					out<=12;
				end
				if(in == 186) begin
					state<=20;
					out<=13;
				end
				if(in == 187) begin
					state<=20;
					out<=14;
				end
				if(in == 188) begin
					state<=20;
					out<=15;
				end
				if(in == 189) begin
					state<=20;
					out<=16;
				end
				if(in == 190) begin
					state<=20;
					out<=17;
				end
				if(in == 191) begin
					state<=20;
					out<=18;
				end
				if(in == 192) begin
					state<=20;
					out<=19;
				end
				if(in == 193) begin
					state<=20;
					out<=20;
				end
				if(in == 194) begin
					state<=20;
					out<=21;
				end
				if(in == 195) begin
					state<=20;
					out<=22;
				end
				if(in == 196) begin
					state<=20;
					out<=23;
				end
				if(in == 197) begin
					state<=20;
					out<=24;
				end
				if(in == 198) begin
					state<=20;
					out<=25;
				end
				if(in == 199) begin
					state<=20;
					out<=26;
				end
				if(in == 200) begin
					state<=20;
					out<=27;
				end
				if(in == 201) begin
					state<=20;
					out<=28;
				end
				if(in == 202) begin
					state<=20;
					out<=29;
				end
				if(in == 203) begin
					state<=20;
					out<=30;
				end
				if(in == 204) begin
					state<=20;
					out<=31;
				end
				if(in == 205) begin
					state<=20;
					out<=32;
				end
				if(in == 206) begin
					state<=20;
					out<=33;
				end
				if(in == 207) begin
					state<=20;
					out<=34;
				end
				if(in == 208) begin
					state<=20;
					out<=35;
				end
				if(in == 209) begin
					state<=20;
					out<=36;
				end
				if(in == 210) begin
					state<=20;
					out<=37;
				end
				if(in == 211) begin
					state<=20;
					out<=38;
				end
				if(in == 212) begin
					state<=20;
					out<=39;
				end
				if(in == 213) begin
					state<=20;
					out<=40;
				end
				if(in == 214) begin
					state<=20;
					out<=41;
				end
				if(in == 215) begin
					state<=20;
					out<=42;
				end
				if(in == 216) begin
					state<=20;
					out<=43;
				end
				if(in == 217) begin
					state<=20;
					out<=44;
				end
				if(in == 218) begin
					state<=20;
					out<=45;
				end
				if(in == 219) begin
					state<=20;
					out<=46;
				end
				if(in == 220) begin
					state<=20;
					out<=47;
				end
				if(in == 221) begin
					state<=2;
					out<=48;
				end
				if(in == 222) begin
					state<=2;
					out<=49;
				end
				if(in == 223) begin
					state<=2;
					out<=50;
				end
				if(in == 224) begin
					state<=2;
					out<=51;
				end
				if(in == 225) begin
					state<=2;
					out<=52;
				end
				if(in == 226) begin
					state<=2;
					out<=53;
				end
				if(in == 227) begin
					state<=2;
					out<=54;
				end
				if(in == 228) begin
					state<=2;
					out<=55;
				end
				if(in == 229) begin
					state<=2;
					out<=56;
				end
				if(in == 230) begin
					state<=2;
					out<=57;
				end
				if(in == 231) begin
					state<=2;
					out<=58;
				end
				if(in == 232) begin
					state<=2;
					out<=59;
				end
				if(in == 233) begin
					state<=3;
					out<=60;
				end
				if(in == 234) begin
					state<=19;
					out<=61;
				end
				if(in == 235) begin
					state<=3;
					out<=62;
				end
				if(in == 236) begin
					state<=20;
					out<=63;
				end
				if(in == 237) begin
					state<=3;
					out<=64;
				end
				if(in == 238) begin
					state<=20;
					out<=65;
				end
				if(in == 239) begin
					state<=20;
					out<=66;
				end
				if(in == 240) begin
					state<=20;
					out<=67;
				end
				if(in == 241) begin
					state<=20;
					out<=68;
				end
				if(in == 242) begin
					state<=20;
					out<=69;
				end
				if(in == 243) begin
					state<=20;
					out<=70;
				end
				if(in == 244) begin
					state<=20;
					out<=71;
				end
				if(in == 245) begin
					state<=20;
					out<=72;
				end
				if(in == 246) begin
					state<=20;
					out<=73;
				end
				if(in == 247) begin
					state<=20;
					out<=74;
				end
				if(in == 248) begin
					state<=20;
					out<=75;
				end
				if(in == 249) begin
					state<=20;
					out<=76;
				end
				if(in == 250) begin
					state<=20;
					out<=77;
				end
				if(in == 251) begin
					state<=20;
					out<=78;
				end
				if(in == 252) begin
					state<=20;
					out<=79;
				end
				if(in == 253) begin
					state<=20;
					out<=80;
				end
				if(in == 254) begin
					state<=20;
					out<=81;
				end
				if(in == 255) begin
					state<=20;
					out<=82;
				end
				if(in == 256) begin
					state<=20;
					out<=83;
				end
				if(in == 257) begin
					state<=20;
					out<=84;
				end
				if(in == 258) begin
					state<=20;
					out<=85;
				end
				if(in == 259) begin
					state<=20;
					out<=86;
				end
				if(in == 260) begin
					state<=20;
					out<=87;
				end
				if(in == 261) begin
					state<=20;
					out<=88;
				end
				if(in == 262) begin
					state<=20;
					out<=89;
				end
				if(in == 263) begin
					state<=20;
					out<=90;
				end
				if(in == 264) begin
					state<=20;
					out<=91;
				end
				if(in == 265) begin
					state<=20;
					out<=92;
				end
				if(in == 266) begin
					state<=20;
					out<=93;
				end
				if(in == 267) begin
					state<=20;
					out<=94;
				end
				if(in == 268) begin
					state<=20;
					out<=95;
				end
				if(in == 269) begin
					state<=20;
					out<=96;
				end
				if(in == 270) begin
					state<=20;
					out<=97;
				end
				if(in == 271) begin
					state<=20;
					out<=98;
				end
				if(in == 272) begin
					state<=20;
					out<=99;
				end
				if(in == 273) begin
					state<=20;
					out<=100;
				end
				if(in == 274) begin
					state<=20;
					out<=101;
				end
				if(in == 275) begin
					state<=20;
					out<=102;
				end
				if(in == 276) begin
					state<=20;
					out<=103;
				end
				if(in == 277) begin
					state<=20;
					out<=104;
				end
				if(in == 278) begin
					state<=20;
					out<=105;
				end
				if(in == 279) begin
					state<=20;
					out<=106;
				end
				if(in == 280) begin
					state<=20;
					out<=107;
				end
				if(in == 281) begin
					state<=20;
					out<=108;
				end
				if(in == 282) begin
					state<=20;
					out<=109;
				end
				if(in == 283) begin
					state<=20;
					out<=110;
				end
				if(in == 284) begin
					state<=20;
					out<=111;
				end
				if(in == 285) begin
					state<=3;
					out<=112;
				end
				if(in == 286) begin
					state<=19;
					out<=113;
				end
				if(in == 287) begin
					state<=3;
					out<=114;
				end
				if(in == 288) begin
					state<=20;
					out<=115;
				end
				if(in == 289) begin
					state<=3;
					out<=116;
				end
				if(in == 290) begin
					state<=20;
					out<=117;
				end
				if(in == 291) begin
					state<=20;
					out<=118;
				end
				if(in == 292) begin
					state<=20;
					out<=119;
				end
				if(in == 293) begin
					state<=20;
					out<=120;
				end
				if(in == 294) begin
					state<=20;
					out<=121;
				end
				if(in == 295) begin
					state<=20;
					out<=122;
				end
				if(in == 296) begin
					state<=20;
					out<=123;
				end
				if(in == 297) begin
					state<=20;
					out<=124;
				end
				if(in == 298) begin
					state<=20;
					out<=125;
				end
				if(in == 299) begin
					state<=20;
					out<=126;
				end
				if(in == 300) begin
					state<=20;
					out<=127;
				end
				if(in == 301) begin
					state<=20;
					out<=128;
				end
				if(in == 302) begin
					state<=20;
					out<=129;
				end
				if(in == 303) begin
					state<=20;
					out<=130;
				end
				if(in == 304) begin
					state<=20;
					out<=131;
				end
				if(in == 305) begin
					state<=20;
					out<=132;
				end
				if(in == 306) begin
					state<=20;
					out<=133;
				end
				if(in == 307) begin
					state<=20;
					out<=134;
				end
				if(in == 308) begin
					state<=20;
					out<=135;
				end
				if(in == 309) begin
					state<=20;
					out<=136;
				end
				if(in == 310) begin
					state<=20;
					out<=137;
				end
				if(in == 311) begin
					state<=20;
					out<=138;
				end
				if(in == 312) begin
					state<=20;
					out<=139;
				end
				if(in == 313) begin
					state<=20;
					out<=140;
				end
				if(in == 314) begin
					state<=20;
					out<=141;
				end
				if(in == 315) begin
					state<=20;
					out<=142;
				end
				if(in == 316) begin
					state<=20;
					out<=143;
				end
				if(in == 317) begin
					state<=20;
					out<=144;
				end
				if(in == 318) begin
					state<=20;
					out<=145;
				end
				if(in == 319) begin
					state<=20;
					out<=146;
				end
				if(in == 320) begin
					state<=20;
					out<=147;
				end
				if(in == 321) begin
					state<=20;
					out<=148;
				end
				if(in == 322) begin
					state<=20;
					out<=149;
				end
				if(in == 323) begin
					state<=20;
					out<=150;
				end
				if(in == 324) begin
					state<=20;
					out<=151;
				end
				if(in == 325) begin
					state<=20;
					out<=152;
				end
				if(in == 326) begin
					state<=20;
					out<=153;
				end
				if(in == 327) begin
					state<=20;
					out<=154;
				end
				if(in == 328) begin
					state<=20;
					out<=155;
				end
				if(in == 329) begin
					state<=20;
					out<=156;
				end
				if(in == 330) begin
					state<=20;
					out<=157;
				end
				if(in == 331) begin
					state<=20;
					out<=158;
				end
				if(in == 332) begin
					state<=20;
					out<=159;
				end
				if(in == 333) begin
					state<=20;
					out<=160;
				end
				if(in == 334) begin
					state<=20;
					out<=161;
				end
				if(in == 335) begin
					state<=20;
					out<=162;
				end
				if(in == 336) begin
					state<=20;
					out<=163;
				end
				if(in == 337) begin
					state<=2;
					out<=164;
				end
				if(in == 338) begin
					state<=2;
					out<=165;
				end
				if(in == 339) begin
					state<=2;
					out<=166;
				end
				if(in == 340) begin
					state<=2;
					out<=167;
				end
				if(in == 341) begin
					state<=2;
					out<=168;
				end
				if(in == 342) begin
					state<=2;
					out<=169;
				end
				if(in == 343) begin
					state<=2;
					out<=170;
				end
				if(in == 344) begin
					state<=2;
					out<=171;
				end
				if(in == 345) begin
					state<=2;
					out<=172;
				end
				if(in == 346) begin
					state<=2;
					out<=173;
				end
				if(in == 347) begin
					state<=2;
					out<=174;
				end
				if(in == 348) begin
					state<=2;
					out<=175;
				end
				if(in == 349) begin
					state<=3;
					out<=176;
				end
				if(in == 350) begin
					state<=19;
					out<=177;
				end
				if(in == 351) begin
					state<=3;
					out<=178;
				end
				if(in == 352) begin
					state<=20;
					out<=179;
				end
				if(in == 353) begin
					state<=3;
					out<=180;
				end
				if(in == 354) begin
					state<=20;
					out<=181;
				end
				if(in == 355) begin
					state<=20;
					out<=182;
				end
				if(in == 356) begin
					state<=20;
					out<=183;
				end
				if(in == 357) begin
					state<=20;
					out<=184;
				end
				if(in == 358) begin
					state<=20;
					out<=185;
				end
				if(in == 359) begin
					state<=20;
					out<=186;
				end
				if(in == 360) begin
					state<=20;
					out<=187;
				end
				if(in == 361) begin
					state<=20;
					out<=188;
				end
				if(in == 362) begin
					state<=20;
					out<=189;
				end
				if(in == 363) begin
					state<=20;
					out<=190;
				end
				if(in == 364) begin
					state<=20;
					out<=191;
				end
				if(in == 365) begin
					state<=20;
					out<=192;
				end
				if(in == 366) begin
					state<=20;
					out<=193;
				end
				if(in == 367) begin
					state<=20;
					out<=194;
				end
				if(in == 368) begin
					state<=20;
					out<=195;
				end
				if(in == 369) begin
					state<=20;
					out<=196;
				end
				if(in == 370) begin
					state<=20;
					out<=197;
				end
				if(in == 371) begin
					state<=20;
					out<=198;
				end
				if(in == 372) begin
					state<=20;
					out<=199;
				end
				if(in == 373) begin
					state<=20;
					out<=200;
				end
				if(in == 374) begin
					state<=20;
					out<=201;
				end
				if(in == 375) begin
					state<=20;
					out<=202;
				end
				if(in == 376) begin
					state<=20;
					out<=203;
				end
				if(in == 377) begin
					state<=20;
					out<=204;
				end
				if(in == 378) begin
					state<=20;
					out<=205;
				end
				if(in == 379) begin
					state<=20;
					out<=206;
				end
				if(in == 380) begin
					state<=20;
					out<=207;
				end
				if(in == 381) begin
					state<=20;
					out<=208;
				end
				if(in == 382) begin
					state<=20;
					out<=209;
				end
				if(in == 383) begin
					state<=20;
					out<=210;
				end
				if(in == 384) begin
					state<=20;
					out<=211;
				end
				if(in == 385) begin
					state<=20;
					out<=212;
				end
				if(in == 386) begin
					state<=20;
					out<=213;
				end
				if(in == 387) begin
					state<=20;
					out<=214;
				end
				if(in == 388) begin
					state<=20;
					out<=215;
				end
				if(in == 389) begin
					state<=20;
					out<=216;
				end
				if(in == 390) begin
					state<=20;
					out<=217;
				end
				if(in == 391) begin
					state<=20;
					out<=218;
				end
				if(in == 392) begin
					state<=20;
					out<=219;
				end
				if(in == 393) begin
					state<=20;
					out<=220;
				end
				if(in == 394) begin
					state<=20;
					out<=221;
				end
				if(in == 395) begin
					state<=20;
					out<=222;
				end
				if(in == 396) begin
					state<=20;
					out<=223;
				end
				if(in == 397) begin
					state<=20;
					out<=224;
				end
				if(in == 398) begin
					state<=20;
					out<=225;
				end
				if(in == 399) begin
					state<=20;
					out<=226;
				end
				if(in == 400) begin
					state<=20;
					out<=227;
				end
				if(in == 401) begin
					state<=3;
					out<=228;
				end
				if(in == 402) begin
					state<=19;
					out<=229;
				end
				if(in == 403) begin
					state<=3;
					out<=230;
				end
				if(in == 404) begin
					state<=20;
					out<=231;
				end
				if(in == 405) begin
					state<=3;
					out<=232;
				end
				if(in == 406) begin
					state<=20;
					out<=233;
				end
				if(in == 407) begin
					state<=20;
					out<=234;
				end
				if(in == 408) begin
					state<=20;
					out<=235;
				end
				if(in == 409) begin
					state<=20;
					out<=236;
				end
				if(in == 410) begin
					state<=20;
					out<=237;
				end
				if(in == 411) begin
					state<=20;
					out<=238;
				end
				if(in == 412) begin
					state<=20;
					out<=239;
				end
				if(in == 413) begin
					state<=20;
					out<=240;
				end
				if(in == 414) begin
					state<=20;
					out<=241;
				end
				if(in == 415) begin
					state<=20;
					out<=242;
				end
				if(in == 416) begin
					state<=20;
					out<=243;
				end
				if(in == 417) begin
					state<=20;
					out<=244;
				end
				if(in == 418) begin
					state<=20;
					out<=245;
				end
				if(in == 419) begin
					state<=20;
					out<=246;
				end
				if(in == 420) begin
					state<=20;
					out<=247;
				end
				if(in == 421) begin
					state<=20;
					out<=248;
				end
				if(in == 422) begin
					state<=20;
					out<=249;
				end
				if(in == 423) begin
					state<=20;
					out<=250;
				end
				if(in == 424) begin
					state<=20;
					out<=251;
				end
				if(in == 425) begin
					state<=20;
					out<=252;
				end
				if(in == 426) begin
					state<=20;
					out<=253;
				end
				if(in == 427) begin
					state<=20;
					out<=254;
				end
				if(in == 428) begin
					state<=20;
					out<=255;
				end
				if(in == 429) begin
					state<=20;
					out<=0;
				end
				if(in == 430) begin
					state<=20;
					out<=1;
				end
				if(in == 431) begin
					state<=20;
					out<=2;
				end
				if(in == 432) begin
					state<=20;
					out<=3;
				end
				if(in == 433) begin
					state<=20;
					out<=4;
				end
				if(in == 434) begin
					state<=20;
					out<=5;
				end
				if(in == 435) begin
					state<=20;
					out<=6;
				end
				if(in == 436) begin
					state<=20;
					out<=7;
				end
				if(in == 437) begin
					state<=20;
					out<=8;
				end
				if(in == 438) begin
					state<=20;
					out<=9;
				end
				if(in == 439) begin
					state<=20;
					out<=10;
				end
				if(in == 440) begin
					state<=20;
					out<=11;
				end
				if(in == 441) begin
					state<=20;
					out<=12;
				end
				if(in == 442) begin
					state<=20;
					out<=13;
				end
				if(in == 443) begin
					state<=20;
					out<=14;
				end
				if(in == 444) begin
					state<=20;
					out<=15;
				end
				if(in == 445) begin
					state<=20;
					out<=16;
				end
				if(in == 446) begin
					state<=20;
					out<=17;
				end
				if(in == 447) begin
					state<=20;
					out<=18;
				end
				if(in == 448) begin
					state<=20;
					out<=19;
				end
				if(in == 449) begin
					state<=20;
					out<=20;
				end
				if(in == 450) begin
					state<=20;
					out<=21;
				end
				if(in == 451) begin
					state<=20;
					out<=22;
				end
				if(in == 452) begin
					state<=20;
					out<=23;
				end
				if(in == 453) begin
					state<=2;
					out<=24;
				end
				if(in == 454) begin
					state<=2;
					out<=25;
				end
				if(in == 455) begin
					state<=2;
					out<=26;
				end
				if(in == 456) begin
					state<=2;
					out<=27;
				end
				if(in == 457) begin
					state<=2;
					out<=28;
				end
				if(in == 458) begin
					state<=2;
					out<=29;
				end
				if(in == 459) begin
					state<=2;
					out<=30;
				end
				if(in == 460) begin
					state<=2;
					out<=31;
				end
				if(in == 461) begin
					state<=2;
					out<=32;
				end
				if(in == 462) begin
					state<=2;
					out<=33;
				end
				if(in == 463) begin
					state<=2;
					out<=34;
				end
				if(in == 464) begin
					state<=2;
					out<=35;
				end
				if(in == 465) begin
					state<=3;
					out<=36;
				end
				if(in == 466) begin
					state<=19;
					out<=37;
				end
				if(in == 467) begin
					state<=3;
					out<=38;
				end
				if(in == 468) begin
					state<=20;
					out<=39;
				end
				if(in == 469) begin
					state<=3;
					out<=40;
				end
				if(in == 470) begin
					state<=20;
					out<=41;
				end
				if(in == 471) begin
					state<=20;
					out<=42;
				end
				if(in == 472) begin
					state<=20;
					out<=43;
				end
				if(in == 473) begin
					state<=20;
					out<=44;
				end
				if(in == 474) begin
					state<=20;
					out<=45;
				end
				if(in == 475) begin
					state<=20;
					out<=46;
				end
				if(in == 476) begin
					state<=20;
					out<=47;
				end
				if(in == 477) begin
					state<=20;
					out<=48;
				end
				if(in == 478) begin
					state<=20;
					out<=49;
				end
				if(in == 479) begin
					state<=20;
					out<=50;
				end
				if(in == 480) begin
					state<=20;
					out<=51;
				end
				if(in == 481) begin
					state<=20;
					out<=52;
				end
				if(in == 482) begin
					state<=20;
					out<=53;
				end
				if(in == 483) begin
					state<=20;
					out<=54;
				end
				if(in == 484) begin
					state<=20;
					out<=55;
				end
				if(in == 485) begin
					state<=20;
					out<=56;
				end
				if(in == 486) begin
					state<=20;
					out<=57;
				end
				if(in == 487) begin
					state<=20;
					out<=58;
				end
				if(in == 488) begin
					state<=20;
					out<=59;
				end
				if(in == 489) begin
					state<=20;
					out<=60;
				end
				if(in == 490) begin
					state<=20;
					out<=61;
				end
				if(in == 491) begin
					state<=20;
					out<=62;
				end
				if(in == 492) begin
					state<=20;
					out<=63;
				end
				if(in == 493) begin
					state<=20;
					out<=64;
				end
				if(in == 494) begin
					state<=20;
					out<=65;
				end
				if(in == 495) begin
					state<=20;
					out<=66;
				end
				if(in == 496) begin
					state<=20;
					out<=67;
				end
				if(in == 497) begin
					state<=20;
					out<=68;
				end
				if(in == 498) begin
					state<=20;
					out<=69;
				end
				if(in == 499) begin
					state<=20;
					out<=70;
				end
				if(in == 500) begin
					state<=20;
					out<=71;
				end
				if(in == 501) begin
					state<=20;
					out<=72;
				end
				if(in == 502) begin
					state<=20;
					out<=73;
				end
				if(in == 503) begin
					state<=20;
					out<=74;
				end
				if(in == 504) begin
					state<=20;
					out<=75;
				end
				if(in == 505) begin
					state<=20;
					out<=76;
				end
				if(in == 506) begin
					state<=20;
					out<=77;
				end
				if(in == 507) begin
					state<=20;
					out<=78;
				end
				if(in == 508) begin
					state<=20;
					out<=79;
				end
				if(in == 509) begin
					state<=20;
					out<=80;
				end
				if(in == 510) begin
					state<=20;
					out<=81;
				end
				if(in == 511) begin
					state<=20;
					out<=82;
				end
				if(in == 512) begin
					state<=20;
					out<=83;
				end
				if(in == 513) begin
					state<=20;
					out<=84;
				end
				if(in == 514) begin
					state<=20;
					out<=85;
				end
				if(in == 515) begin
					state<=20;
					out<=86;
				end
				if(in == 516) begin
					state<=20;
					out<=87;
				end
				if(in == 517) begin
					state<=3;
					out<=88;
				end
				if(in == 518) begin
					state<=19;
					out<=89;
				end
				if(in == 519) begin
					state<=3;
					out<=90;
				end
				if(in == 520) begin
					state<=20;
					out<=91;
				end
				if(in == 521) begin
					state<=3;
					out<=92;
				end
				if(in == 522) begin
					state<=20;
					out<=93;
				end
				if(in == 523) begin
					state<=20;
					out<=94;
				end
				if(in == 524) begin
					state<=20;
					out<=95;
				end
				if(in == 525) begin
					state<=20;
					out<=96;
				end
				if(in == 526) begin
					state<=20;
					out<=97;
				end
				if(in == 527) begin
					state<=20;
					out<=98;
				end
				if(in == 528) begin
					state<=20;
					out<=99;
				end
				if(in == 529) begin
					state<=20;
					out<=100;
				end
				if(in == 530) begin
					state<=20;
					out<=101;
				end
				if(in == 531) begin
					state<=20;
					out<=102;
				end
				if(in == 532) begin
					state<=20;
					out<=103;
				end
				if(in == 533) begin
					state<=20;
					out<=104;
				end
				if(in == 534) begin
					state<=20;
					out<=105;
				end
				if(in == 535) begin
					state<=20;
					out<=106;
				end
				if(in == 536) begin
					state<=20;
					out<=107;
				end
				if(in == 537) begin
					state<=20;
					out<=108;
				end
				if(in == 538) begin
					state<=20;
					out<=109;
				end
				if(in == 539) begin
					state<=20;
					out<=110;
				end
				if(in == 540) begin
					state<=20;
					out<=111;
				end
				if(in == 541) begin
					state<=20;
					out<=112;
				end
				if(in == 542) begin
					state<=20;
					out<=113;
				end
				if(in == 543) begin
					state<=20;
					out<=114;
				end
				if(in == 544) begin
					state<=20;
					out<=115;
				end
				if(in == 545) begin
					state<=20;
					out<=116;
				end
				if(in == 546) begin
					state<=20;
					out<=117;
				end
				if(in == 547) begin
					state<=20;
					out<=118;
				end
				if(in == 548) begin
					state<=20;
					out<=119;
				end
				if(in == 549) begin
					state<=20;
					out<=120;
				end
				if(in == 550) begin
					state<=20;
					out<=121;
				end
				if(in == 551) begin
					state<=20;
					out<=122;
				end
				if(in == 552) begin
					state<=20;
					out<=123;
				end
				if(in == 553) begin
					state<=20;
					out<=124;
				end
				if(in == 554) begin
					state<=20;
					out<=125;
				end
				if(in == 555) begin
					state<=20;
					out<=126;
				end
				if(in == 556) begin
					state<=20;
					out<=127;
				end
				if(in == 557) begin
					state<=20;
					out<=128;
				end
				if(in == 558) begin
					state<=20;
					out<=129;
				end
				if(in == 559) begin
					state<=20;
					out<=130;
				end
				if(in == 560) begin
					state<=20;
					out<=131;
				end
				if(in == 561) begin
					state<=20;
					out<=132;
				end
				if(in == 562) begin
					state<=20;
					out<=133;
				end
				if(in == 563) begin
					state<=20;
					out<=134;
				end
				if(in == 564) begin
					state<=20;
					out<=135;
				end
				if(in == 565) begin
					state<=20;
					out<=136;
				end
				if(in == 566) begin
					state<=20;
					out<=137;
				end
				if(in == 567) begin
					state<=20;
					out<=138;
				end
				if(in == 568) begin
					state<=20;
					out<=139;
				end
				if(in == 569) begin
					state<=2;
					out<=140;
				end
				if(in == 570) begin
					state<=2;
					out<=141;
				end
				if(in == 571) begin
					state<=2;
					out<=142;
				end
				if(in == 572) begin
					state<=2;
					out<=143;
				end
				if(in == 573) begin
					state<=2;
					out<=144;
				end
				if(in == 574) begin
					state<=2;
					out<=145;
				end
				if(in == 575) begin
					state<=2;
					out<=146;
				end
				if(in == 576) begin
					state<=2;
					out<=147;
				end
				if(in == 577) begin
					state<=2;
					out<=148;
				end
				if(in == 578) begin
					state<=2;
					out<=149;
				end
				if(in == 579) begin
					state<=2;
					out<=150;
				end
				if(in == 580) begin
					state<=2;
					out<=151;
				end
				if(in == 581) begin
					state<=3;
					out<=152;
				end
				if(in == 582) begin
					state<=19;
					out<=153;
				end
				if(in == 583) begin
					state<=3;
					out<=154;
				end
				if(in == 584) begin
					state<=20;
					out<=155;
				end
				if(in == 585) begin
					state<=3;
					out<=156;
				end
				if(in == 586) begin
					state<=20;
					out<=157;
				end
				if(in == 587) begin
					state<=20;
					out<=158;
				end
				if(in == 588) begin
					state<=20;
					out<=159;
				end
				if(in == 589) begin
					state<=20;
					out<=160;
				end
				if(in == 590) begin
					state<=20;
					out<=161;
				end
				if(in == 591) begin
					state<=20;
					out<=162;
				end
				if(in == 592) begin
					state<=20;
					out<=163;
				end
				if(in == 593) begin
					state<=20;
					out<=164;
				end
				if(in == 594) begin
					state<=20;
					out<=165;
				end
				if(in == 595) begin
					state<=20;
					out<=166;
				end
				if(in == 596) begin
					state<=20;
					out<=167;
				end
				if(in == 597) begin
					state<=20;
					out<=168;
				end
				if(in == 598) begin
					state<=20;
					out<=169;
				end
				if(in == 599) begin
					state<=20;
					out<=170;
				end
				if(in == 600) begin
					state<=20;
					out<=171;
				end
				if(in == 601) begin
					state<=20;
					out<=172;
				end
				if(in == 602) begin
					state<=20;
					out<=173;
				end
				if(in == 603) begin
					state<=20;
					out<=174;
				end
				if(in == 604) begin
					state<=20;
					out<=175;
				end
				if(in == 605) begin
					state<=20;
					out<=176;
				end
				if(in == 606) begin
					state<=20;
					out<=177;
				end
				if(in == 607) begin
					state<=20;
					out<=178;
				end
				if(in == 608) begin
					state<=20;
					out<=179;
				end
				if(in == 609) begin
					state<=20;
					out<=180;
				end
				if(in == 610) begin
					state<=20;
					out<=181;
				end
				if(in == 611) begin
					state<=20;
					out<=182;
				end
				if(in == 612) begin
					state<=20;
					out<=183;
				end
				if(in == 613) begin
					state<=20;
					out<=184;
				end
				if(in == 614) begin
					state<=20;
					out<=185;
				end
				if(in == 615) begin
					state<=20;
					out<=186;
				end
				if(in == 616) begin
					state<=20;
					out<=187;
				end
				if(in == 617) begin
					state<=20;
					out<=188;
				end
				if(in == 618) begin
					state<=20;
					out<=189;
				end
				if(in == 619) begin
					state<=20;
					out<=190;
				end
				if(in == 620) begin
					state<=20;
					out<=191;
				end
				if(in == 621) begin
					state<=20;
					out<=192;
				end
				if(in == 622) begin
					state<=20;
					out<=193;
				end
				if(in == 623) begin
					state<=20;
					out<=194;
				end
				if(in == 624) begin
					state<=20;
					out<=195;
				end
				if(in == 625) begin
					state<=20;
					out<=196;
				end
				if(in == 626) begin
					state<=20;
					out<=197;
				end
				if(in == 627) begin
					state<=20;
					out<=198;
				end
				if(in == 628) begin
					state<=20;
					out<=199;
				end
				if(in == 629) begin
					state<=20;
					out<=200;
				end
				if(in == 630) begin
					state<=20;
					out<=201;
				end
				if(in == 631) begin
					state<=20;
					out<=202;
				end
				if(in == 632) begin
					state<=20;
					out<=203;
				end
				if(in == 633) begin
					state<=3;
					out<=204;
				end
				if(in == 634) begin
					state<=19;
					out<=205;
				end
				if(in == 635) begin
					state<=3;
					out<=206;
				end
				if(in == 636) begin
					state<=20;
					out<=207;
				end
				if(in == 637) begin
					state<=3;
					out<=208;
				end
				if(in == 638) begin
					state<=20;
					out<=209;
				end
				if(in == 639) begin
					state<=20;
					out<=210;
				end
				if(in == 640) begin
					state<=20;
					out<=211;
				end
				if(in == 641) begin
					state<=20;
					out<=212;
				end
				if(in == 642) begin
					state<=20;
					out<=213;
				end
				if(in == 643) begin
					state<=20;
					out<=214;
				end
				if(in == 644) begin
					state<=20;
					out<=215;
				end
				if(in == 645) begin
					state<=20;
					out<=216;
				end
				if(in == 646) begin
					state<=20;
					out<=217;
				end
				if(in == 647) begin
					state<=20;
					out<=218;
				end
				if(in == 648) begin
					state<=20;
					out<=219;
				end
				if(in == 649) begin
					state<=20;
					out<=220;
				end
				if(in == 650) begin
					state<=20;
					out<=221;
				end
				if(in == 651) begin
					state<=20;
					out<=222;
				end
				if(in == 652) begin
					state<=20;
					out<=223;
				end
				if(in == 653) begin
					state<=20;
					out<=224;
				end
				if(in == 654) begin
					state<=20;
					out<=225;
				end
				if(in == 655) begin
					state<=20;
					out<=226;
				end
				if(in == 656) begin
					state<=20;
					out<=227;
				end
				if(in == 657) begin
					state<=20;
					out<=228;
				end
				if(in == 658) begin
					state<=20;
					out<=229;
				end
				if(in == 659) begin
					state<=20;
					out<=230;
				end
				if(in == 660) begin
					state<=20;
					out<=231;
				end
				if(in == 661) begin
					state<=20;
					out<=232;
				end
				if(in == 662) begin
					state<=20;
					out<=233;
				end
				if(in == 663) begin
					state<=20;
					out<=234;
				end
				if(in == 664) begin
					state<=20;
					out<=235;
				end
				if(in == 665) begin
					state<=20;
					out<=236;
				end
				if(in == 666) begin
					state<=20;
					out<=237;
				end
				if(in == 667) begin
					state<=20;
					out<=238;
				end
				if(in == 668) begin
					state<=20;
					out<=239;
				end
				if(in == 669) begin
					state<=20;
					out<=240;
				end
				if(in == 670) begin
					state<=20;
					out<=241;
				end
				if(in == 671) begin
					state<=20;
					out<=242;
				end
				if(in == 672) begin
					state<=20;
					out<=243;
				end
				if(in == 673) begin
					state<=20;
					out<=244;
				end
				if(in == 674) begin
					state<=20;
					out<=245;
				end
				if(in == 675) begin
					state<=20;
					out<=246;
				end
				if(in == 676) begin
					state<=20;
					out<=247;
				end
				if(in == 677) begin
					state<=20;
					out<=248;
				end
				if(in == 678) begin
					state<=20;
					out<=249;
				end
				if(in == 679) begin
					state<=20;
					out<=250;
				end
				if(in == 680) begin
					state<=20;
					out<=251;
				end
				if(in == 681) begin
					state<=20;
					out<=252;
				end
				if(in == 682) begin
					state<=20;
					out<=253;
				end
				if(in == 683) begin
					state<=20;
					out<=254;
				end
				if(in == 684) begin
					state<=20;
					out<=255;
				end
				if(in == 685) begin
					state<=2;
					out<=0;
				end
				if(in == 686) begin
					state<=2;
					out<=1;
				end
				if(in == 687) begin
					state<=2;
					out<=2;
				end
				if(in == 688) begin
					state<=2;
					out<=3;
				end
				if(in == 689) begin
					state<=2;
					out<=4;
				end
				if(in == 690) begin
					state<=2;
					out<=5;
				end
				if(in == 691) begin
					state<=2;
					out<=6;
				end
				if(in == 692) begin
					state<=2;
					out<=7;
				end
				if(in == 693) begin
					state<=2;
					out<=8;
				end
				if(in == 694) begin
					state<=2;
					out<=9;
				end
				if(in == 695) begin
					state<=2;
					out<=10;
				end
				if(in == 696) begin
					state<=2;
					out<=11;
				end
				if(in == 697) begin
					state<=3;
					out<=12;
				end
				if(in == 698) begin
					state<=19;
					out<=13;
				end
				if(in == 699) begin
					state<=3;
					out<=14;
				end
				if(in == 700) begin
					state<=20;
					out<=15;
				end
				if(in == 701) begin
					state<=3;
					out<=16;
				end
				if(in == 702) begin
					state<=20;
					out<=17;
				end
				if(in == 703) begin
					state<=20;
					out<=18;
				end
				if(in == 704) begin
					state<=20;
					out<=19;
				end
				if(in == 705) begin
					state<=20;
					out<=20;
				end
				if(in == 706) begin
					state<=20;
					out<=21;
				end
				if(in == 707) begin
					state<=20;
					out<=22;
				end
				if(in == 708) begin
					state<=20;
					out<=23;
				end
				if(in == 709) begin
					state<=20;
					out<=24;
				end
				if(in == 710) begin
					state<=20;
					out<=25;
				end
				if(in == 711) begin
					state<=20;
					out<=26;
				end
				if(in == 712) begin
					state<=20;
					out<=27;
				end
				if(in == 713) begin
					state<=20;
					out<=28;
				end
				if(in == 714) begin
					state<=20;
					out<=29;
				end
				if(in == 715) begin
					state<=20;
					out<=30;
				end
				if(in == 716) begin
					state<=20;
					out<=31;
				end
				if(in == 717) begin
					state<=20;
					out<=32;
				end
				if(in == 718) begin
					state<=20;
					out<=33;
				end
				if(in == 719) begin
					state<=20;
					out<=34;
				end
				if(in == 720) begin
					state<=20;
					out<=35;
				end
				if(in == 721) begin
					state<=20;
					out<=36;
				end
				if(in == 722) begin
					state<=20;
					out<=37;
				end
				if(in == 723) begin
					state<=20;
					out<=38;
				end
				if(in == 724) begin
					state<=20;
					out<=39;
				end
				if(in == 725) begin
					state<=20;
					out<=40;
				end
				if(in == 726) begin
					state<=20;
					out<=41;
				end
				if(in == 727) begin
					state<=20;
					out<=42;
				end
				if(in == 728) begin
					state<=20;
					out<=43;
				end
				if(in == 729) begin
					state<=20;
					out<=44;
				end
				if(in == 730) begin
					state<=20;
					out<=45;
				end
				if(in == 731) begin
					state<=20;
					out<=46;
				end
				if(in == 732) begin
					state<=20;
					out<=47;
				end
				if(in == 733) begin
					state<=20;
					out<=48;
				end
				if(in == 734) begin
					state<=20;
					out<=49;
				end
				if(in == 735) begin
					state<=20;
					out<=50;
				end
				if(in == 736) begin
					state<=20;
					out<=51;
				end
				if(in == 737) begin
					state<=20;
					out<=52;
				end
				if(in == 738) begin
					state<=20;
					out<=53;
				end
				if(in == 739) begin
					state<=20;
					out<=54;
				end
				if(in == 740) begin
					state<=20;
					out<=55;
				end
				if(in == 741) begin
					state<=20;
					out<=56;
				end
				if(in == 742) begin
					state<=20;
					out<=57;
				end
				if(in == 743) begin
					state<=20;
					out<=58;
				end
				if(in == 744) begin
					state<=20;
					out<=59;
				end
				if(in == 745) begin
					state<=20;
					out<=60;
				end
				if(in == 746) begin
					state<=20;
					out<=61;
				end
				if(in == 747) begin
					state<=20;
					out<=62;
				end
				if(in == 748) begin
					state<=20;
					out<=63;
				end
				if(in == 749) begin
					state<=3;
					out<=64;
				end
				if(in == 750) begin
					state<=19;
					out<=65;
				end
				if(in == 751) begin
					state<=3;
					out<=66;
				end
				if(in == 752) begin
					state<=20;
					out<=67;
				end
				if(in == 753) begin
					state<=3;
					out<=68;
				end
				if(in == 754) begin
					state<=20;
					out<=69;
				end
				if(in == 755) begin
					state<=20;
					out<=70;
				end
				if(in == 756) begin
					state<=20;
					out<=71;
				end
				if(in == 757) begin
					state<=20;
					out<=72;
				end
				if(in == 758) begin
					state<=20;
					out<=73;
				end
				if(in == 759) begin
					state<=20;
					out<=74;
				end
				if(in == 760) begin
					state<=20;
					out<=75;
				end
				if(in == 761) begin
					state<=20;
					out<=76;
				end
				if(in == 762) begin
					state<=20;
					out<=77;
				end
				if(in == 763) begin
					state<=20;
					out<=78;
				end
				if(in == 764) begin
					state<=20;
					out<=79;
				end
				if(in == 765) begin
					state<=20;
					out<=80;
				end
				if(in == 766) begin
					state<=20;
					out<=81;
				end
				if(in == 767) begin
					state<=20;
					out<=82;
				end
				if(in == 768) begin
					state<=20;
					out<=83;
				end
				if(in == 769) begin
					state<=20;
					out<=84;
				end
				if(in == 770) begin
					state<=20;
					out<=85;
				end
				if(in == 771) begin
					state<=20;
					out<=86;
				end
				if(in == 772) begin
					state<=20;
					out<=87;
				end
				if(in == 773) begin
					state<=20;
					out<=88;
				end
				if(in == 774) begin
					state<=20;
					out<=89;
				end
				if(in == 775) begin
					state<=20;
					out<=90;
				end
				if(in == 776) begin
					state<=20;
					out<=91;
				end
				if(in == 777) begin
					state<=20;
					out<=92;
				end
				if(in == 778) begin
					state<=20;
					out<=93;
				end
				if(in == 779) begin
					state<=20;
					out<=94;
				end
				if(in == 780) begin
					state<=20;
					out<=95;
				end
				if(in == 781) begin
					state<=20;
					out<=96;
				end
				if(in == 782) begin
					state<=20;
					out<=97;
				end
				if(in == 783) begin
					state<=20;
					out<=98;
				end
				if(in == 784) begin
					state<=20;
					out<=99;
				end
				if(in == 785) begin
					state<=20;
					out<=100;
				end
				if(in == 786) begin
					state<=20;
					out<=101;
				end
				if(in == 787) begin
					state<=20;
					out<=102;
				end
				if(in == 788) begin
					state<=20;
					out<=103;
				end
				if(in == 789) begin
					state<=20;
					out<=104;
				end
				if(in == 790) begin
					state<=20;
					out<=105;
				end
				if(in == 791) begin
					state<=20;
					out<=106;
				end
				if(in == 792) begin
					state<=20;
					out<=107;
				end
				if(in == 793) begin
					state<=20;
					out<=108;
				end
				if(in == 794) begin
					state<=20;
					out<=109;
				end
				if(in == 795) begin
					state<=20;
					out<=110;
				end
				if(in == 796) begin
					state<=20;
					out<=111;
				end
				if(in == 797) begin
					state<=20;
					out<=112;
				end
				if(in == 798) begin
					state<=20;
					out<=113;
				end
				if(in == 799) begin
					state<=20;
					out<=114;
				end
				if(in == 800) begin
					state<=20;
					out<=115;
				end
				if(in == 801) begin
					state<=2;
					out<=116;
				end
				if(in == 802) begin
					state<=2;
					out<=117;
				end
				if(in == 803) begin
					state<=2;
					out<=118;
				end
				if(in == 804) begin
					state<=2;
					out<=119;
				end
				if(in == 805) begin
					state<=2;
					out<=120;
				end
				if(in == 806) begin
					state<=2;
					out<=121;
				end
				if(in == 807) begin
					state<=2;
					out<=122;
				end
				if(in == 808) begin
					state<=2;
					out<=123;
				end
				if(in == 809) begin
					state<=2;
					out<=124;
				end
				if(in == 810) begin
					state<=2;
					out<=125;
				end
				if(in == 811) begin
					state<=2;
					out<=126;
				end
				if(in == 812) begin
					state<=2;
					out<=127;
				end
				if(in == 813) begin
					state<=3;
					out<=128;
				end
				if(in == 814) begin
					state<=19;
					out<=129;
				end
				if(in == 815) begin
					state<=3;
					out<=130;
				end
				if(in == 816) begin
					state<=20;
					out<=131;
				end
				if(in == 817) begin
					state<=3;
					out<=132;
				end
				if(in == 818) begin
					state<=20;
					out<=133;
				end
				if(in == 819) begin
					state<=20;
					out<=134;
				end
				if(in == 820) begin
					state<=20;
					out<=135;
				end
				if(in == 821) begin
					state<=20;
					out<=136;
				end
				if(in == 822) begin
					state<=20;
					out<=137;
				end
				if(in == 823) begin
					state<=20;
					out<=138;
				end
				if(in == 824) begin
					state<=20;
					out<=139;
				end
				if(in == 825) begin
					state<=20;
					out<=140;
				end
				if(in == 826) begin
					state<=20;
					out<=141;
				end
				if(in == 827) begin
					state<=20;
					out<=142;
				end
				if(in == 828) begin
					state<=20;
					out<=143;
				end
				if(in == 829) begin
					state<=20;
					out<=144;
				end
				if(in == 830) begin
					state<=20;
					out<=145;
				end
				if(in == 831) begin
					state<=20;
					out<=146;
				end
				if(in == 832) begin
					state<=20;
					out<=147;
				end
				if(in == 833) begin
					state<=20;
					out<=148;
				end
				if(in == 834) begin
					state<=20;
					out<=149;
				end
				if(in == 835) begin
					state<=20;
					out<=150;
				end
				if(in == 836) begin
					state<=20;
					out<=151;
				end
				if(in == 837) begin
					state<=20;
					out<=152;
				end
				if(in == 838) begin
					state<=20;
					out<=153;
				end
				if(in == 839) begin
					state<=20;
					out<=154;
				end
				if(in == 840) begin
					state<=20;
					out<=155;
				end
				if(in == 841) begin
					state<=20;
					out<=156;
				end
				if(in == 842) begin
					state<=20;
					out<=157;
				end
				if(in == 843) begin
					state<=20;
					out<=158;
				end
				if(in == 844) begin
					state<=20;
					out<=159;
				end
				if(in == 845) begin
					state<=20;
					out<=160;
				end
				if(in == 846) begin
					state<=20;
					out<=161;
				end
				if(in == 847) begin
					state<=20;
					out<=162;
				end
				if(in == 848) begin
					state<=20;
					out<=163;
				end
				if(in == 849) begin
					state<=20;
					out<=164;
				end
				if(in == 850) begin
					state<=20;
					out<=165;
				end
				if(in == 851) begin
					state<=20;
					out<=166;
				end
				if(in == 852) begin
					state<=20;
					out<=167;
				end
				if(in == 853) begin
					state<=20;
					out<=168;
				end
				if(in == 854) begin
					state<=20;
					out<=169;
				end
				if(in == 855) begin
					state<=20;
					out<=170;
				end
				if(in == 856) begin
					state<=20;
					out<=171;
				end
				if(in == 857) begin
					state<=20;
					out<=172;
				end
				if(in == 858) begin
					state<=20;
					out<=173;
				end
				if(in == 859) begin
					state<=20;
					out<=174;
				end
				if(in == 860) begin
					state<=20;
					out<=175;
				end
				if(in == 861) begin
					state<=20;
					out<=176;
				end
				if(in == 862) begin
					state<=20;
					out<=177;
				end
				if(in == 863) begin
					state<=20;
					out<=178;
				end
				if(in == 864) begin
					state<=20;
					out<=179;
				end
				if(in == 865) begin
					state<=3;
					out<=180;
				end
				if(in == 866) begin
					state<=19;
					out<=181;
				end
				if(in == 867) begin
					state<=3;
					out<=182;
				end
				if(in == 868) begin
					state<=20;
					out<=183;
				end
				if(in == 869) begin
					state<=3;
					out<=184;
				end
				if(in == 870) begin
					state<=20;
					out<=185;
				end
				if(in == 871) begin
					state<=20;
					out<=186;
				end
				if(in == 872) begin
					state<=20;
					out<=187;
				end
				if(in == 873) begin
					state<=20;
					out<=188;
				end
				if(in == 874) begin
					state<=20;
					out<=189;
				end
				if(in == 875) begin
					state<=20;
					out<=190;
				end
				if(in == 876) begin
					state<=20;
					out<=191;
				end
				if(in == 877) begin
					state<=20;
					out<=192;
				end
				if(in == 878) begin
					state<=20;
					out<=193;
				end
				if(in == 879) begin
					state<=20;
					out<=194;
				end
				if(in == 880) begin
					state<=20;
					out<=195;
				end
				if(in == 881) begin
					state<=20;
					out<=196;
				end
				if(in == 882) begin
					state<=20;
					out<=197;
				end
				if(in == 883) begin
					state<=20;
					out<=198;
				end
				if(in == 884) begin
					state<=20;
					out<=199;
				end
				if(in == 885) begin
					state<=20;
					out<=200;
				end
				if(in == 886) begin
					state<=20;
					out<=201;
				end
				if(in == 887) begin
					state<=20;
					out<=202;
				end
				if(in == 888) begin
					state<=20;
					out<=203;
				end
				if(in == 889) begin
					state<=20;
					out<=204;
				end
				if(in == 890) begin
					state<=20;
					out<=205;
				end
				if(in == 891) begin
					state<=20;
					out<=206;
				end
				if(in == 892) begin
					state<=20;
					out<=207;
				end
				if(in == 893) begin
					state<=20;
					out<=208;
				end
				if(in == 894) begin
					state<=20;
					out<=209;
				end
				if(in == 895) begin
					state<=20;
					out<=210;
				end
				if(in == 896) begin
					state<=20;
					out<=211;
				end
				if(in == 897) begin
					state<=20;
					out<=212;
				end
				if(in == 898) begin
					state<=20;
					out<=213;
				end
				if(in == 899) begin
					state<=20;
					out<=214;
				end
				if(in == 900) begin
					state<=20;
					out<=215;
				end
				if(in == 901) begin
					state<=20;
					out<=216;
				end
				if(in == 902) begin
					state<=20;
					out<=217;
				end
				if(in == 903) begin
					state<=20;
					out<=218;
				end
				if(in == 904) begin
					state<=20;
					out<=219;
				end
				if(in == 905) begin
					state<=20;
					out<=220;
				end
				if(in == 906) begin
					state<=20;
					out<=221;
				end
				if(in == 907) begin
					state<=20;
					out<=222;
				end
				if(in == 908) begin
					state<=20;
					out<=223;
				end
				if(in == 909) begin
					state<=20;
					out<=224;
				end
				if(in == 910) begin
					state<=20;
					out<=225;
				end
				if(in == 911) begin
					state<=20;
					out<=226;
				end
				if(in == 912) begin
					state<=20;
					out<=227;
				end
				if(in == 913) begin
					state<=20;
					out<=228;
				end
				if(in == 914) begin
					state<=20;
					out<=229;
				end
				if(in == 915) begin
					state<=20;
					out<=230;
				end
				if(in == 916) begin
					state<=20;
					out<=231;
				end
				if(in == 917) begin
					state<=2;
					out<=232;
				end
				if(in == 918) begin
					state<=2;
					out<=233;
				end
				if(in == 919) begin
					state<=2;
					out<=234;
				end
				if(in == 920) begin
					state<=2;
					out<=235;
				end
				if(in == 921) begin
					state<=2;
					out<=236;
				end
				if(in == 922) begin
					state<=2;
					out<=237;
				end
				if(in == 923) begin
					state<=2;
					out<=238;
				end
				if(in == 924) begin
					state<=2;
					out<=239;
				end
				if(in == 925) begin
					state<=2;
					out<=240;
				end
				if(in == 926) begin
					state<=2;
					out<=241;
				end
				if(in == 927) begin
					state<=2;
					out<=242;
				end
				if(in == 928) begin
					state<=2;
					out<=243;
				end
			end
			20: begin
				if(in == 0) begin
					state<=3;
					out<=244;
				end
				if(in == 1) begin
					state<=1;
					out<=245;
				end
				if(in == 2) begin
					state<=20;
					out<=246;
				end
				if(in == 3) begin
					state<=3;
					out<=247;
				end
				if(in == 4) begin
					state<=21;
					out<=248;
				end
				if(in == 5) begin
					state<=3;
					out<=249;
				end
				if(in == 6) begin
					state<=21;
					out<=250;
				end
				if(in == 7) begin
					state<=21;
					out<=251;
				end
				if(in == 8) begin
					state<=21;
					out<=252;
				end
				if(in == 9) begin
					state<=21;
					out<=253;
				end
				if(in == 10) begin
					state<=21;
					out<=254;
				end
				if(in == 11) begin
					state<=21;
					out<=255;
				end
				if(in == 12) begin
					state<=21;
					out<=0;
				end
				if(in == 13) begin
					state<=21;
					out<=1;
				end
				if(in == 14) begin
					state<=21;
					out<=2;
				end
				if(in == 15) begin
					state<=21;
					out<=3;
				end
				if(in == 16) begin
					state<=21;
					out<=4;
				end
				if(in == 17) begin
					state<=21;
					out<=5;
				end
				if(in == 18) begin
					state<=21;
					out<=6;
				end
				if(in == 19) begin
					state<=21;
					out<=7;
				end
				if(in == 20) begin
					state<=21;
					out<=8;
				end
				if(in == 21) begin
					state<=21;
					out<=9;
				end
				if(in == 22) begin
					state<=21;
					out<=10;
				end
				if(in == 23) begin
					state<=21;
					out<=11;
				end
				if(in == 24) begin
					state<=21;
					out<=12;
				end
				if(in == 25) begin
					state<=21;
					out<=13;
				end
				if(in == 26) begin
					state<=21;
					out<=14;
				end
				if(in == 27) begin
					state<=21;
					out<=15;
				end
				if(in == 28) begin
					state<=21;
					out<=16;
				end
				if(in == 29) begin
					state<=21;
					out<=17;
				end
				if(in == 30) begin
					state<=21;
					out<=18;
				end
				if(in == 31) begin
					state<=21;
					out<=19;
				end
				if(in == 32) begin
					state<=21;
					out<=20;
				end
				if(in == 33) begin
					state<=21;
					out<=21;
				end
				if(in == 34) begin
					state<=21;
					out<=22;
				end
				if(in == 35) begin
					state<=21;
					out<=23;
				end
				if(in == 36) begin
					state<=21;
					out<=24;
				end
				if(in == 37) begin
					state<=21;
					out<=25;
				end
				if(in == 38) begin
					state<=21;
					out<=26;
				end
				if(in == 39) begin
					state<=21;
					out<=27;
				end
				if(in == 40) begin
					state<=21;
					out<=28;
				end
				if(in == 41) begin
					state<=21;
					out<=29;
				end
				if(in == 42) begin
					state<=21;
					out<=30;
				end
				if(in == 43) begin
					state<=21;
					out<=31;
				end
				if(in == 44) begin
					state<=21;
					out<=32;
				end
				if(in == 45) begin
					state<=21;
					out<=33;
				end
				if(in == 46) begin
					state<=21;
					out<=34;
				end
				if(in == 47) begin
					state<=21;
					out<=35;
				end
				if(in == 48) begin
					state<=21;
					out<=36;
				end
				if(in == 49) begin
					state<=21;
					out<=37;
				end
				if(in == 50) begin
					state<=21;
					out<=38;
				end
				if(in == 51) begin
					state<=21;
					out<=39;
				end
				if(in == 52) begin
					state<=21;
					out<=40;
				end
				if(in == 53) begin
					state<=3;
					out<=41;
				end
				if(in == 54) begin
					state<=20;
					out<=42;
				end
				if(in == 55) begin
					state<=3;
					out<=43;
				end
				if(in == 56) begin
					state<=21;
					out<=44;
				end
				if(in == 57) begin
					state<=3;
					out<=45;
				end
				if(in == 58) begin
					state<=21;
					out<=46;
				end
				if(in == 59) begin
					state<=21;
					out<=47;
				end
				if(in == 60) begin
					state<=21;
					out<=48;
				end
				if(in == 61) begin
					state<=21;
					out<=49;
				end
				if(in == 62) begin
					state<=21;
					out<=50;
				end
				if(in == 63) begin
					state<=21;
					out<=51;
				end
				if(in == 64) begin
					state<=21;
					out<=52;
				end
				if(in == 65) begin
					state<=21;
					out<=53;
				end
				if(in == 66) begin
					state<=21;
					out<=54;
				end
				if(in == 67) begin
					state<=21;
					out<=55;
				end
				if(in == 68) begin
					state<=21;
					out<=56;
				end
				if(in == 69) begin
					state<=21;
					out<=57;
				end
				if(in == 70) begin
					state<=21;
					out<=58;
				end
				if(in == 71) begin
					state<=21;
					out<=59;
				end
				if(in == 72) begin
					state<=21;
					out<=60;
				end
				if(in == 73) begin
					state<=21;
					out<=61;
				end
				if(in == 74) begin
					state<=21;
					out<=62;
				end
				if(in == 75) begin
					state<=21;
					out<=63;
				end
				if(in == 76) begin
					state<=21;
					out<=64;
				end
				if(in == 77) begin
					state<=21;
					out<=65;
				end
				if(in == 78) begin
					state<=21;
					out<=66;
				end
				if(in == 79) begin
					state<=21;
					out<=67;
				end
				if(in == 80) begin
					state<=21;
					out<=68;
				end
				if(in == 81) begin
					state<=21;
					out<=69;
				end
				if(in == 82) begin
					state<=21;
					out<=70;
				end
				if(in == 83) begin
					state<=21;
					out<=71;
				end
				if(in == 84) begin
					state<=21;
					out<=72;
				end
				if(in == 85) begin
					state<=21;
					out<=73;
				end
				if(in == 86) begin
					state<=21;
					out<=74;
				end
				if(in == 87) begin
					state<=21;
					out<=75;
				end
				if(in == 88) begin
					state<=21;
					out<=76;
				end
				if(in == 89) begin
					state<=21;
					out<=77;
				end
				if(in == 90) begin
					state<=21;
					out<=78;
				end
				if(in == 91) begin
					state<=21;
					out<=79;
				end
				if(in == 92) begin
					state<=21;
					out<=80;
				end
				if(in == 93) begin
					state<=21;
					out<=81;
				end
				if(in == 94) begin
					state<=21;
					out<=82;
				end
				if(in == 95) begin
					state<=21;
					out<=83;
				end
				if(in == 96) begin
					state<=21;
					out<=84;
				end
				if(in == 97) begin
					state<=21;
					out<=85;
				end
				if(in == 98) begin
					state<=21;
					out<=86;
				end
				if(in == 99) begin
					state<=21;
					out<=87;
				end
				if(in == 100) begin
					state<=21;
					out<=88;
				end
				if(in == 101) begin
					state<=21;
					out<=89;
				end
				if(in == 102) begin
					state<=21;
					out<=90;
				end
				if(in == 103) begin
					state<=21;
					out<=91;
				end
				if(in == 104) begin
					state<=21;
					out<=92;
				end
				if(in == 105) begin
					state<=2;
					out<=93;
				end
				if(in == 106) begin
					state<=2;
					out<=94;
				end
				if(in == 107) begin
					state<=2;
					out<=95;
				end
				if(in == 108) begin
					state<=2;
					out<=96;
				end
				if(in == 109) begin
					state<=2;
					out<=97;
				end
				if(in == 110) begin
					state<=2;
					out<=98;
				end
				if(in == 111) begin
					state<=2;
					out<=99;
				end
				if(in == 112) begin
					state<=2;
					out<=100;
				end
				if(in == 113) begin
					state<=2;
					out<=101;
				end
				if(in == 114) begin
					state<=2;
					out<=102;
				end
				if(in == 115) begin
					state<=2;
					out<=103;
				end
				if(in == 116) begin
					state<=2;
					out<=104;
				end
				if(in == 117) begin
					state<=3;
					out<=105;
				end
				if(in == 118) begin
					state<=20;
					out<=106;
				end
				if(in == 119) begin
					state<=3;
					out<=107;
				end
				if(in == 120) begin
					state<=21;
					out<=108;
				end
				if(in == 121) begin
					state<=3;
					out<=109;
				end
				if(in == 122) begin
					state<=21;
					out<=110;
				end
				if(in == 123) begin
					state<=21;
					out<=111;
				end
				if(in == 124) begin
					state<=21;
					out<=112;
				end
				if(in == 125) begin
					state<=21;
					out<=113;
				end
				if(in == 126) begin
					state<=21;
					out<=114;
				end
				if(in == 127) begin
					state<=21;
					out<=115;
				end
				if(in == 128) begin
					state<=21;
					out<=116;
				end
				if(in == 129) begin
					state<=21;
					out<=117;
				end
				if(in == 130) begin
					state<=21;
					out<=118;
				end
				if(in == 131) begin
					state<=21;
					out<=119;
				end
				if(in == 132) begin
					state<=21;
					out<=120;
				end
				if(in == 133) begin
					state<=21;
					out<=121;
				end
				if(in == 134) begin
					state<=21;
					out<=122;
				end
				if(in == 135) begin
					state<=21;
					out<=123;
				end
				if(in == 136) begin
					state<=21;
					out<=124;
				end
				if(in == 137) begin
					state<=21;
					out<=125;
				end
				if(in == 138) begin
					state<=21;
					out<=126;
				end
				if(in == 139) begin
					state<=21;
					out<=127;
				end
				if(in == 140) begin
					state<=21;
					out<=128;
				end
				if(in == 141) begin
					state<=21;
					out<=129;
				end
				if(in == 142) begin
					state<=21;
					out<=130;
				end
				if(in == 143) begin
					state<=21;
					out<=131;
				end
				if(in == 144) begin
					state<=21;
					out<=132;
				end
				if(in == 145) begin
					state<=21;
					out<=133;
				end
				if(in == 146) begin
					state<=21;
					out<=134;
				end
				if(in == 147) begin
					state<=21;
					out<=135;
				end
				if(in == 148) begin
					state<=21;
					out<=136;
				end
				if(in == 149) begin
					state<=21;
					out<=137;
				end
				if(in == 150) begin
					state<=21;
					out<=138;
				end
				if(in == 151) begin
					state<=21;
					out<=139;
				end
				if(in == 152) begin
					state<=21;
					out<=140;
				end
				if(in == 153) begin
					state<=21;
					out<=141;
				end
				if(in == 154) begin
					state<=21;
					out<=142;
				end
				if(in == 155) begin
					state<=21;
					out<=143;
				end
				if(in == 156) begin
					state<=21;
					out<=144;
				end
				if(in == 157) begin
					state<=21;
					out<=145;
				end
				if(in == 158) begin
					state<=21;
					out<=146;
				end
				if(in == 159) begin
					state<=21;
					out<=147;
				end
				if(in == 160) begin
					state<=21;
					out<=148;
				end
				if(in == 161) begin
					state<=21;
					out<=149;
				end
				if(in == 162) begin
					state<=21;
					out<=150;
				end
				if(in == 163) begin
					state<=21;
					out<=151;
				end
				if(in == 164) begin
					state<=21;
					out<=152;
				end
				if(in == 165) begin
					state<=21;
					out<=153;
				end
				if(in == 166) begin
					state<=21;
					out<=154;
				end
				if(in == 167) begin
					state<=21;
					out<=155;
				end
				if(in == 168) begin
					state<=21;
					out<=156;
				end
				if(in == 169) begin
					state<=3;
					out<=157;
				end
				if(in == 170) begin
					state<=20;
					out<=158;
				end
				if(in == 171) begin
					state<=3;
					out<=159;
				end
				if(in == 172) begin
					state<=21;
					out<=160;
				end
				if(in == 173) begin
					state<=3;
					out<=161;
				end
				if(in == 174) begin
					state<=21;
					out<=162;
				end
				if(in == 175) begin
					state<=21;
					out<=163;
				end
				if(in == 176) begin
					state<=21;
					out<=164;
				end
				if(in == 177) begin
					state<=21;
					out<=165;
				end
				if(in == 178) begin
					state<=21;
					out<=166;
				end
				if(in == 179) begin
					state<=21;
					out<=167;
				end
				if(in == 180) begin
					state<=21;
					out<=168;
				end
				if(in == 181) begin
					state<=21;
					out<=169;
				end
				if(in == 182) begin
					state<=21;
					out<=170;
				end
				if(in == 183) begin
					state<=21;
					out<=171;
				end
				if(in == 184) begin
					state<=21;
					out<=172;
				end
				if(in == 185) begin
					state<=21;
					out<=173;
				end
				if(in == 186) begin
					state<=21;
					out<=174;
				end
				if(in == 187) begin
					state<=21;
					out<=175;
				end
				if(in == 188) begin
					state<=21;
					out<=176;
				end
				if(in == 189) begin
					state<=21;
					out<=177;
				end
				if(in == 190) begin
					state<=21;
					out<=178;
				end
				if(in == 191) begin
					state<=21;
					out<=179;
				end
				if(in == 192) begin
					state<=21;
					out<=180;
				end
				if(in == 193) begin
					state<=21;
					out<=181;
				end
				if(in == 194) begin
					state<=21;
					out<=182;
				end
				if(in == 195) begin
					state<=21;
					out<=183;
				end
				if(in == 196) begin
					state<=21;
					out<=184;
				end
				if(in == 197) begin
					state<=21;
					out<=185;
				end
				if(in == 198) begin
					state<=21;
					out<=186;
				end
				if(in == 199) begin
					state<=21;
					out<=187;
				end
				if(in == 200) begin
					state<=21;
					out<=188;
				end
				if(in == 201) begin
					state<=21;
					out<=189;
				end
				if(in == 202) begin
					state<=21;
					out<=190;
				end
				if(in == 203) begin
					state<=21;
					out<=191;
				end
				if(in == 204) begin
					state<=21;
					out<=192;
				end
				if(in == 205) begin
					state<=21;
					out<=193;
				end
				if(in == 206) begin
					state<=21;
					out<=194;
				end
				if(in == 207) begin
					state<=21;
					out<=195;
				end
				if(in == 208) begin
					state<=21;
					out<=196;
				end
				if(in == 209) begin
					state<=21;
					out<=197;
				end
				if(in == 210) begin
					state<=21;
					out<=198;
				end
				if(in == 211) begin
					state<=21;
					out<=199;
				end
				if(in == 212) begin
					state<=21;
					out<=200;
				end
				if(in == 213) begin
					state<=21;
					out<=201;
				end
				if(in == 214) begin
					state<=21;
					out<=202;
				end
				if(in == 215) begin
					state<=21;
					out<=203;
				end
				if(in == 216) begin
					state<=21;
					out<=204;
				end
				if(in == 217) begin
					state<=21;
					out<=205;
				end
				if(in == 218) begin
					state<=21;
					out<=206;
				end
				if(in == 219) begin
					state<=21;
					out<=207;
				end
				if(in == 220) begin
					state<=21;
					out<=208;
				end
				if(in == 221) begin
					state<=2;
					out<=209;
				end
				if(in == 222) begin
					state<=2;
					out<=210;
				end
				if(in == 223) begin
					state<=2;
					out<=211;
				end
				if(in == 224) begin
					state<=2;
					out<=212;
				end
				if(in == 225) begin
					state<=2;
					out<=213;
				end
				if(in == 226) begin
					state<=2;
					out<=214;
				end
				if(in == 227) begin
					state<=2;
					out<=215;
				end
				if(in == 228) begin
					state<=2;
					out<=216;
				end
				if(in == 229) begin
					state<=2;
					out<=217;
				end
				if(in == 230) begin
					state<=2;
					out<=218;
				end
				if(in == 231) begin
					state<=2;
					out<=219;
				end
				if(in == 232) begin
					state<=2;
					out<=220;
				end
				if(in == 233) begin
					state<=3;
					out<=221;
				end
				if(in == 234) begin
					state<=20;
					out<=222;
				end
				if(in == 235) begin
					state<=3;
					out<=223;
				end
				if(in == 236) begin
					state<=21;
					out<=224;
				end
				if(in == 237) begin
					state<=3;
					out<=225;
				end
				if(in == 238) begin
					state<=21;
					out<=226;
				end
				if(in == 239) begin
					state<=21;
					out<=227;
				end
				if(in == 240) begin
					state<=21;
					out<=228;
				end
				if(in == 241) begin
					state<=21;
					out<=229;
				end
				if(in == 242) begin
					state<=21;
					out<=230;
				end
				if(in == 243) begin
					state<=21;
					out<=231;
				end
				if(in == 244) begin
					state<=21;
					out<=232;
				end
				if(in == 245) begin
					state<=21;
					out<=233;
				end
				if(in == 246) begin
					state<=21;
					out<=234;
				end
				if(in == 247) begin
					state<=21;
					out<=235;
				end
				if(in == 248) begin
					state<=21;
					out<=236;
				end
				if(in == 249) begin
					state<=21;
					out<=237;
				end
				if(in == 250) begin
					state<=21;
					out<=238;
				end
				if(in == 251) begin
					state<=21;
					out<=239;
				end
				if(in == 252) begin
					state<=21;
					out<=240;
				end
				if(in == 253) begin
					state<=21;
					out<=241;
				end
				if(in == 254) begin
					state<=21;
					out<=242;
				end
				if(in == 255) begin
					state<=21;
					out<=243;
				end
				if(in == 256) begin
					state<=21;
					out<=244;
				end
				if(in == 257) begin
					state<=21;
					out<=245;
				end
				if(in == 258) begin
					state<=21;
					out<=246;
				end
				if(in == 259) begin
					state<=21;
					out<=247;
				end
				if(in == 260) begin
					state<=21;
					out<=248;
				end
				if(in == 261) begin
					state<=21;
					out<=249;
				end
				if(in == 262) begin
					state<=21;
					out<=250;
				end
				if(in == 263) begin
					state<=21;
					out<=251;
				end
				if(in == 264) begin
					state<=21;
					out<=252;
				end
				if(in == 265) begin
					state<=21;
					out<=253;
				end
				if(in == 266) begin
					state<=21;
					out<=254;
				end
				if(in == 267) begin
					state<=21;
					out<=255;
				end
				if(in == 268) begin
					state<=21;
					out<=0;
				end
				if(in == 269) begin
					state<=21;
					out<=1;
				end
				if(in == 270) begin
					state<=21;
					out<=2;
				end
				if(in == 271) begin
					state<=21;
					out<=3;
				end
				if(in == 272) begin
					state<=21;
					out<=4;
				end
				if(in == 273) begin
					state<=21;
					out<=5;
				end
				if(in == 274) begin
					state<=21;
					out<=6;
				end
				if(in == 275) begin
					state<=21;
					out<=7;
				end
				if(in == 276) begin
					state<=21;
					out<=8;
				end
				if(in == 277) begin
					state<=21;
					out<=9;
				end
				if(in == 278) begin
					state<=21;
					out<=10;
				end
				if(in == 279) begin
					state<=21;
					out<=11;
				end
				if(in == 280) begin
					state<=21;
					out<=12;
				end
				if(in == 281) begin
					state<=21;
					out<=13;
				end
				if(in == 282) begin
					state<=21;
					out<=14;
				end
				if(in == 283) begin
					state<=21;
					out<=15;
				end
				if(in == 284) begin
					state<=21;
					out<=16;
				end
				if(in == 285) begin
					state<=3;
					out<=17;
				end
				if(in == 286) begin
					state<=20;
					out<=18;
				end
				if(in == 287) begin
					state<=3;
					out<=19;
				end
				if(in == 288) begin
					state<=21;
					out<=20;
				end
				if(in == 289) begin
					state<=3;
					out<=21;
				end
				if(in == 290) begin
					state<=21;
					out<=22;
				end
				if(in == 291) begin
					state<=21;
					out<=23;
				end
				if(in == 292) begin
					state<=21;
					out<=24;
				end
				if(in == 293) begin
					state<=21;
					out<=25;
				end
				if(in == 294) begin
					state<=21;
					out<=26;
				end
				if(in == 295) begin
					state<=21;
					out<=27;
				end
				if(in == 296) begin
					state<=21;
					out<=28;
				end
				if(in == 297) begin
					state<=21;
					out<=29;
				end
				if(in == 298) begin
					state<=21;
					out<=30;
				end
				if(in == 299) begin
					state<=21;
					out<=31;
				end
				if(in == 300) begin
					state<=21;
					out<=32;
				end
				if(in == 301) begin
					state<=21;
					out<=33;
				end
				if(in == 302) begin
					state<=21;
					out<=34;
				end
				if(in == 303) begin
					state<=21;
					out<=35;
				end
				if(in == 304) begin
					state<=21;
					out<=36;
				end
				if(in == 305) begin
					state<=21;
					out<=37;
				end
				if(in == 306) begin
					state<=21;
					out<=38;
				end
				if(in == 307) begin
					state<=21;
					out<=39;
				end
				if(in == 308) begin
					state<=21;
					out<=40;
				end
				if(in == 309) begin
					state<=21;
					out<=41;
				end
				if(in == 310) begin
					state<=21;
					out<=42;
				end
				if(in == 311) begin
					state<=21;
					out<=43;
				end
				if(in == 312) begin
					state<=21;
					out<=44;
				end
				if(in == 313) begin
					state<=21;
					out<=45;
				end
				if(in == 314) begin
					state<=21;
					out<=46;
				end
				if(in == 315) begin
					state<=21;
					out<=47;
				end
				if(in == 316) begin
					state<=21;
					out<=48;
				end
				if(in == 317) begin
					state<=21;
					out<=49;
				end
				if(in == 318) begin
					state<=21;
					out<=50;
				end
				if(in == 319) begin
					state<=21;
					out<=51;
				end
				if(in == 320) begin
					state<=21;
					out<=52;
				end
				if(in == 321) begin
					state<=21;
					out<=53;
				end
				if(in == 322) begin
					state<=21;
					out<=54;
				end
				if(in == 323) begin
					state<=21;
					out<=55;
				end
				if(in == 324) begin
					state<=21;
					out<=56;
				end
				if(in == 325) begin
					state<=21;
					out<=57;
				end
				if(in == 326) begin
					state<=21;
					out<=58;
				end
				if(in == 327) begin
					state<=21;
					out<=59;
				end
				if(in == 328) begin
					state<=21;
					out<=60;
				end
				if(in == 329) begin
					state<=21;
					out<=61;
				end
				if(in == 330) begin
					state<=21;
					out<=62;
				end
				if(in == 331) begin
					state<=21;
					out<=63;
				end
				if(in == 332) begin
					state<=21;
					out<=64;
				end
				if(in == 333) begin
					state<=21;
					out<=65;
				end
				if(in == 334) begin
					state<=21;
					out<=66;
				end
				if(in == 335) begin
					state<=21;
					out<=67;
				end
				if(in == 336) begin
					state<=21;
					out<=68;
				end
				if(in == 337) begin
					state<=2;
					out<=69;
				end
				if(in == 338) begin
					state<=2;
					out<=70;
				end
				if(in == 339) begin
					state<=2;
					out<=71;
				end
				if(in == 340) begin
					state<=2;
					out<=72;
				end
				if(in == 341) begin
					state<=2;
					out<=73;
				end
				if(in == 342) begin
					state<=2;
					out<=74;
				end
				if(in == 343) begin
					state<=2;
					out<=75;
				end
				if(in == 344) begin
					state<=2;
					out<=76;
				end
				if(in == 345) begin
					state<=2;
					out<=77;
				end
				if(in == 346) begin
					state<=2;
					out<=78;
				end
				if(in == 347) begin
					state<=2;
					out<=79;
				end
				if(in == 348) begin
					state<=2;
					out<=80;
				end
				if(in == 349) begin
					state<=3;
					out<=81;
				end
				if(in == 350) begin
					state<=20;
					out<=82;
				end
				if(in == 351) begin
					state<=3;
					out<=83;
				end
				if(in == 352) begin
					state<=21;
					out<=84;
				end
				if(in == 353) begin
					state<=3;
					out<=85;
				end
				if(in == 354) begin
					state<=21;
					out<=86;
				end
				if(in == 355) begin
					state<=21;
					out<=87;
				end
				if(in == 356) begin
					state<=21;
					out<=88;
				end
				if(in == 357) begin
					state<=21;
					out<=89;
				end
				if(in == 358) begin
					state<=21;
					out<=90;
				end
				if(in == 359) begin
					state<=21;
					out<=91;
				end
				if(in == 360) begin
					state<=21;
					out<=92;
				end
				if(in == 361) begin
					state<=21;
					out<=93;
				end
				if(in == 362) begin
					state<=21;
					out<=94;
				end
				if(in == 363) begin
					state<=21;
					out<=95;
				end
				if(in == 364) begin
					state<=21;
					out<=96;
				end
				if(in == 365) begin
					state<=21;
					out<=97;
				end
				if(in == 366) begin
					state<=21;
					out<=98;
				end
				if(in == 367) begin
					state<=21;
					out<=99;
				end
				if(in == 368) begin
					state<=21;
					out<=100;
				end
				if(in == 369) begin
					state<=21;
					out<=101;
				end
				if(in == 370) begin
					state<=21;
					out<=102;
				end
				if(in == 371) begin
					state<=21;
					out<=103;
				end
				if(in == 372) begin
					state<=21;
					out<=104;
				end
				if(in == 373) begin
					state<=21;
					out<=105;
				end
				if(in == 374) begin
					state<=21;
					out<=106;
				end
				if(in == 375) begin
					state<=21;
					out<=107;
				end
				if(in == 376) begin
					state<=21;
					out<=108;
				end
				if(in == 377) begin
					state<=21;
					out<=109;
				end
				if(in == 378) begin
					state<=21;
					out<=110;
				end
				if(in == 379) begin
					state<=21;
					out<=111;
				end
				if(in == 380) begin
					state<=21;
					out<=112;
				end
				if(in == 381) begin
					state<=21;
					out<=113;
				end
				if(in == 382) begin
					state<=21;
					out<=114;
				end
				if(in == 383) begin
					state<=21;
					out<=115;
				end
				if(in == 384) begin
					state<=21;
					out<=116;
				end
				if(in == 385) begin
					state<=21;
					out<=117;
				end
				if(in == 386) begin
					state<=21;
					out<=118;
				end
				if(in == 387) begin
					state<=21;
					out<=119;
				end
				if(in == 388) begin
					state<=21;
					out<=120;
				end
				if(in == 389) begin
					state<=21;
					out<=121;
				end
				if(in == 390) begin
					state<=21;
					out<=122;
				end
				if(in == 391) begin
					state<=21;
					out<=123;
				end
				if(in == 392) begin
					state<=21;
					out<=124;
				end
				if(in == 393) begin
					state<=21;
					out<=125;
				end
				if(in == 394) begin
					state<=21;
					out<=126;
				end
				if(in == 395) begin
					state<=21;
					out<=127;
				end
				if(in == 396) begin
					state<=21;
					out<=128;
				end
				if(in == 397) begin
					state<=21;
					out<=129;
				end
				if(in == 398) begin
					state<=21;
					out<=130;
				end
				if(in == 399) begin
					state<=21;
					out<=131;
				end
				if(in == 400) begin
					state<=21;
					out<=132;
				end
				if(in == 401) begin
					state<=3;
					out<=133;
				end
				if(in == 402) begin
					state<=20;
					out<=134;
				end
				if(in == 403) begin
					state<=3;
					out<=135;
				end
				if(in == 404) begin
					state<=21;
					out<=136;
				end
				if(in == 405) begin
					state<=3;
					out<=137;
				end
				if(in == 406) begin
					state<=21;
					out<=138;
				end
				if(in == 407) begin
					state<=21;
					out<=139;
				end
				if(in == 408) begin
					state<=21;
					out<=140;
				end
				if(in == 409) begin
					state<=21;
					out<=141;
				end
				if(in == 410) begin
					state<=21;
					out<=142;
				end
				if(in == 411) begin
					state<=21;
					out<=143;
				end
				if(in == 412) begin
					state<=21;
					out<=144;
				end
				if(in == 413) begin
					state<=21;
					out<=145;
				end
				if(in == 414) begin
					state<=21;
					out<=146;
				end
				if(in == 415) begin
					state<=21;
					out<=147;
				end
				if(in == 416) begin
					state<=21;
					out<=148;
				end
				if(in == 417) begin
					state<=21;
					out<=149;
				end
				if(in == 418) begin
					state<=21;
					out<=150;
				end
				if(in == 419) begin
					state<=21;
					out<=151;
				end
				if(in == 420) begin
					state<=21;
					out<=152;
				end
				if(in == 421) begin
					state<=21;
					out<=153;
				end
				if(in == 422) begin
					state<=21;
					out<=154;
				end
				if(in == 423) begin
					state<=21;
					out<=155;
				end
				if(in == 424) begin
					state<=21;
					out<=156;
				end
				if(in == 425) begin
					state<=21;
					out<=157;
				end
				if(in == 426) begin
					state<=21;
					out<=158;
				end
				if(in == 427) begin
					state<=21;
					out<=159;
				end
				if(in == 428) begin
					state<=21;
					out<=160;
				end
				if(in == 429) begin
					state<=21;
					out<=161;
				end
				if(in == 430) begin
					state<=21;
					out<=162;
				end
				if(in == 431) begin
					state<=21;
					out<=163;
				end
				if(in == 432) begin
					state<=21;
					out<=164;
				end
				if(in == 433) begin
					state<=21;
					out<=165;
				end
				if(in == 434) begin
					state<=21;
					out<=166;
				end
				if(in == 435) begin
					state<=21;
					out<=167;
				end
				if(in == 436) begin
					state<=21;
					out<=168;
				end
				if(in == 437) begin
					state<=21;
					out<=169;
				end
				if(in == 438) begin
					state<=21;
					out<=170;
				end
				if(in == 439) begin
					state<=21;
					out<=171;
				end
				if(in == 440) begin
					state<=21;
					out<=172;
				end
				if(in == 441) begin
					state<=21;
					out<=173;
				end
				if(in == 442) begin
					state<=21;
					out<=174;
				end
				if(in == 443) begin
					state<=21;
					out<=175;
				end
				if(in == 444) begin
					state<=21;
					out<=176;
				end
				if(in == 445) begin
					state<=21;
					out<=177;
				end
				if(in == 446) begin
					state<=21;
					out<=178;
				end
				if(in == 447) begin
					state<=21;
					out<=179;
				end
				if(in == 448) begin
					state<=21;
					out<=180;
				end
				if(in == 449) begin
					state<=21;
					out<=181;
				end
				if(in == 450) begin
					state<=21;
					out<=182;
				end
				if(in == 451) begin
					state<=21;
					out<=183;
				end
				if(in == 452) begin
					state<=21;
					out<=184;
				end
				if(in == 453) begin
					state<=2;
					out<=185;
				end
				if(in == 454) begin
					state<=2;
					out<=186;
				end
				if(in == 455) begin
					state<=2;
					out<=187;
				end
				if(in == 456) begin
					state<=2;
					out<=188;
				end
				if(in == 457) begin
					state<=2;
					out<=189;
				end
				if(in == 458) begin
					state<=2;
					out<=190;
				end
				if(in == 459) begin
					state<=2;
					out<=191;
				end
				if(in == 460) begin
					state<=2;
					out<=192;
				end
				if(in == 461) begin
					state<=2;
					out<=193;
				end
				if(in == 462) begin
					state<=2;
					out<=194;
				end
				if(in == 463) begin
					state<=2;
					out<=195;
				end
				if(in == 464) begin
					state<=2;
					out<=196;
				end
				if(in == 465) begin
					state<=3;
					out<=197;
				end
				if(in == 466) begin
					state<=20;
					out<=198;
				end
				if(in == 467) begin
					state<=3;
					out<=199;
				end
				if(in == 468) begin
					state<=21;
					out<=200;
				end
				if(in == 469) begin
					state<=3;
					out<=201;
				end
				if(in == 470) begin
					state<=21;
					out<=202;
				end
				if(in == 471) begin
					state<=21;
					out<=203;
				end
				if(in == 472) begin
					state<=21;
					out<=204;
				end
				if(in == 473) begin
					state<=21;
					out<=205;
				end
				if(in == 474) begin
					state<=21;
					out<=206;
				end
				if(in == 475) begin
					state<=21;
					out<=207;
				end
				if(in == 476) begin
					state<=21;
					out<=208;
				end
				if(in == 477) begin
					state<=21;
					out<=209;
				end
				if(in == 478) begin
					state<=21;
					out<=210;
				end
				if(in == 479) begin
					state<=21;
					out<=211;
				end
				if(in == 480) begin
					state<=21;
					out<=212;
				end
				if(in == 481) begin
					state<=21;
					out<=213;
				end
				if(in == 482) begin
					state<=21;
					out<=214;
				end
				if(in == 483) begin
					state<=21;
					out<=215;
				end
				if(in == 484) begin
					state<=21;
					out<=216;
				end
				if(in == 485) begin
					state<=21;
					out<=217;
				end
				if(in == 486) begin
					state<=21;
					out<=218;
				end
				if(in == 487) begin
					state<=21;
					out<=219;
				end
				if(in == 488) begin
					state<=21;
					out<=220;
				end
				if(in == 489) begin
					state<=21;
					out<=221;
				end
				if(in == 490) begin
					state<=21;
					out<=222;
				end
				if(in == 491) begin
					state<=21;
					out<=223;
				end
				if(in == 492) begin
					state<=21;
					out<=224;
				end
				if(in == 493) begin
					state<=21;
					out<=225;
				end
				if(in == 494) begin
					state<=21;
					out<=226;
				end
				if(in == 495) begin
					state<=21;
					out<=227;
				end
				if(in == 496) begin
					state<=21;
					out<=228;
				end
				if(in == 497) begin
					state<=21;
					out<=229;
				end
				if(in == 498) begin
					state<=21;
					out<=230;
				end
				if(in == 499) begin
					state<=21;
					out<=231;
				end
				if(in == 500) begin
					state<=21;
					out<=232;
				end
				if(in == 501) begin
					state<=21;
					out<=233;
				end
				if(in == 502) begin
					state<=21;
					out<=234;
				end
				if(in == 503) begin
					state<=21;
					out<=235;
				end
				if(in == 504) begin
					state<=21;
					out<=236;
				end
				if(in == 505) begin
					state<=21;
					out<=237;
				end
				if(in == 506) begin
					state<=21;
					out<=238;
				end
				if(in == 507) begin
					state<=21;
					out<=239;
				end
				if(in == 508) begin
					state<=21;
					out<=240;
				end
				if(in == 509) begin
					state<=21;
					out<=241;
				end
				if(in == 510) begin
					state<=21;
					out<=242;
				end
				if(in == 511) begin
					state<=21;
					out<=243;
				end
				if(in == 512) begin
					state<=21;
					out<=244;
				end
				if(in == 513) begin
					state<=21;
					out<=245;
				end
				if(in == 514) begin
					state<=21;
					out<=246;
				end
				if(in == 515) begin
					state<=21;
					out<=247;
				end
				if(in == 516) begin
					state<=21;
					out<=248;
				end
				if(in == 517) begin
					state<=3;
					out<=249;
				end
				if(in == 518) begin
					state<=20;
					out<=250;
				end
				if(in == 519) begin
					state<=3;
					out<=251;
				end
				if(in == 520) begin
					state<=21;
					out<=252;
				end
				if(in == 521) begin
					state<=3;
					out<=253;
				end
				if(in == 522) begin
					state<=21;
					out<=254;
				end
				if(in == 523) begin
					state<=21;
					out<=255;
				end
				if(in == 524) begin
					state<=21;
					out<=0;
				end
				if(in == 525) begin
					state<=21;
					out<=1;
				end
				if(in == 526) begin
					state<=21;
					out<=2;
				end
				if(in == 527) begin
					state<=21;
					out<=3;
				end
				if(in == 528) begin
					state<=21;
					out<=4;
				end
				if(in == 529) begin
					state<=21;
					out<=5;
				end
				if(in == 530) begin
					state<=21;
					out<=6;
				end
				if(in == 531) begin
					state<=21;
					out<=7;
				end
				if(in == 532) begin
					state<=21;
					out<=8;
				end
				if(in == 533) begin
					state<=21;
					out<=9;
				end
				if(in == 534) begin
					state<=21;
					out<=10;
				end
				if(in == 535) begin
					state<=21;
					out<=11;
				end
				if(in == 536) begin
					state<=21;
					out<=12;
				end
				if(in == 537) begin
					state<=21;
					out<=13;
				end
				if(in == 538) begin
					state<=21;
					out<=14;
				end
				if(in == 539) begin
					state<=21;
					out<=15;
				end
				if(in == 540) begin
					state<=21;
					out<=16;
				end
				if(in == 541) begin
					state<=21;
					out<=17;
				end
				if(in == 542) begin
					state<=21;
					out<=18;
				end
				if(in == 543) begin
					state<=21;
					out<=19;
				end
				if(in == 544) begin
					state<=21;
					out<=20;
				end
				if(in == 545) begin
					state<=21;
					out<=21;
				end
				if(in == 546) begin
					state<=21;
					out<=22;
				end
				if(in == 547) begin
					state<=21;
					out<=23;
				end
				if(in == 548) begin
					state<=21;
					out<=24;
				end
				if(in == 549) begin
					state<=21;
					out<=25;
				end
				if(in == 550) begin
					state<=21;
					out<=26;
				end
				if(in == 551) begin
					state<=21;
					out<=27;
				end
				if(in == 552) begin
					state<=21;
					out<=28;
				end
				if(in == 553) begin
					state<=21;
					out<=29;
				end
				if(in == 554) begin
					state<=21;
					out<=30;
				end
				if(in == 555) begin
					state<=21;
					out<=31;
				end
				if(in == 556) begin
					state<=21;
					out<=32;
				end
				if(in == 557) begin
					state<=21;
					out<=33;
				end
				if(in == 558) begin
					state<=21;
					out<=34;
				end
				if(in == 559) begin
					state<=21;
					out<=35;
				end
				if(in == 560) begin
					state<=21;
					out<=36;
				end
				if(in == 561) begin
					state<=21;
					out<=37;
				end
				if(in == 562) begin
					state<=21;
					out<=38;
				end
				if(in == 563) begin
					state<=21;
					out<=39;
				end
				if(in == 564) begin
					state<=21;
					out<=40;
				end
				if(in == 565) begin
					state<=21;
					out<=41;
				end
				if(in == 566) begin
					state<=21;
					out<=42;
				end
				if(in == 567) begin
					state<=21;
					out<=43;
				end
				if(in == 568) begin
					state<=21;
					out<=44;
				end
				if(in == 569) begin
					state<=2;
					out<=45;
				end
				if(in == 570) begin
					state<=2;
					out<=46;
				end
				if(in == 571) begin
					state<=2;
					out<=47;
				end
				if(in == 572) begin
					state<=2;
					out<=48;
				end
				if(in == 573) begin
					state<=2;
					out<=49;
				end
				if(in == 574) begin
					state<=2;
					out<=50;
				end
				if(in == 575) begin
					state<=2;
					out<=51;
				end
				if(in == 576) begin
					state<=2;
					out<=52;
				end
				if(in == 577) begin
					state<=2;
					out<=53;
				end
				if(in == 578) begin
					state<=2;
					out<=54;
				end
				if(in == 579) begin
					state<=2;
					out<=55;
				end
				if(in == 580) begin
					state<=2;
					out<=56;
				end
				if(in == 581) begin
					state<=3;
					out<=57;
				end
				if(in == 582) begin
					state<=20;
					out<=58;
				end
				if(in == 583) begin
					state<=3;
					out<=59;
				end
				if(in == 584) begin
					state<=21;
					out<=60;
				end
				if(in == 585) begin
					state<=3;
					out<=61;
				end
				if(in == 586) begin
					state<=21;
					out<=62;
				end
				if(in == 587) begin
					state<=21;
					out<=63;
				end
				if(in == 588) begin
					state<=21;
					out<=64;
				end
				if(in == 589) begin
					state<=21;
					out<=65;
				end
				if(in == 590) begin
					state<=21;
					out<=66;
				end
				if(in == 591) begin
					state<=21;
					out<=67;
				end
				if(in == 592) begin
					state<=21;
					out<=68;
				end
				if(in == 593) begin
					state<=21;
					out<=69;
				end
				if(in == 594) begin
					state<=21;
					out<=70;
				end
				if(in == 595) begin
					state<=21;
					out<=71;
				end
				if(in == 596) begin
					state<=21;
					out<=72;
				end
				if(in == 597) begin
					state<=21;
					out<=73;
				end
				if(in == 598) begin
					state<=21;
					out<=74;
				end
				if(in == 599) begin
					state<=21;
					out<=75;
				end
				if(in == 600) begin
					state<=21;
					out<=76;
				end
				if(in == 601) begin
					state<=21;
					out<=77;
				end
				if(in == 602) begin
					state<=21;
					out<=78;
				end
				if(in == 603) begin
					state<=21;
					out<=79;
				end
				if(in == 604) begin
					state<=21;
					out<=80;
				end
				if(in == 605) begin
					state<=21;
					out<=81;
				end
				if(in == 606) begin
					state<=21;
					out<=82;
				end
				if(in == 607) begin
					state<=21;
					out<=83;
				end
				if(in == 608) begin
					state<=21;
					out<=84;
				end
				if(in == 609) begin
					state<=21;
					out<=85;
				end
				if(in == 610) begin
					state<=21;
					out<=86;
				end
				if(in == 611) begin
					state<=21;
					out<=87;
				end
				if(in == 612) begin
					state<=21;
					out<=88;
				end
				if(in == 613) begin
					state<=21;
					out<=89;
				end
				if(in == 614) begin
					state<=21;
					out<=90;
				end
				if(in == 615) begin
					state<=21;
					out<=91;
				end
				if(in == 616) begin
					state<=21;
					out<=92;
				end
				if(in == 617) begin
					state<=21;
					out<=93;
				end
				if(in == 618) begin
					state<=21;
					out<=94;
				end
				if(in == 619) begin
					state<=21;
					out<=95;
				end
				if(in == 620) begin
					state<=21;
					out<=96;
				end
				if(in == 621) begin
					state<=21;
					out<=97;
				end
				if(in == 622) begin
					state<=21;
					out<=98;
				end
				if(in == 623) begin
					state<=21;
					out<=99;
				end
				if(in == 624) begin
					state<=21;
					out<=100;
				end
				if(in == 625) begin
					state<=21;
					out<=101;
				end
				if(in == 626) begin
					state<=21;
					out<=102;
				end
				if(in == 627) begin
					state<=21;
					out<=103;
				end
				if(in == 628) begin
					state<=21;
					out<=104;
				end
				if(in == 629) begin
					state<=21;
					out<=105;
				end
				if(in == 630) begin
					state<=21;
					out<=106;
				end
				if(in == 631) begin
					state<=21;
					out<=107;
				end
				if(in == 632) begin
					state<=21;
					out<=108;
				end
				if(in == 633) begin
					state<=3;
					out<=109;
				end
				if(in == 634) begin
					state<=20;
					out<=110;
				end
				if(in == 635) begin
					state<=3;
					out<=111;
				end
				if(in == 636) begin
					state<=21;
					out<=112;
				end
				if(in == 637) begin
					state<=3;
					out<=113;
				end
				if(in == 638) begin
					state<=21;
					out<=114;
				end
				if(in == 639) begin
					state<=21;
					out<=115;
				end
				if(in == 640) begin
					state<=21;
					out<=116;
				end
				if(in == 641) begin
					state<=21;
					out<=117;
				end
				if(in == 642) begin
					state<=21;
					out<=118;
				end
				if(in == 643) begin
					state<=21;
					out<=119;
				end
				if(in == 644) begin
					state<=21;
					out<=120;
				end
				if(in == 645) begin
					state<=21;
					out<=121;
				end
				if(in == 646) begin
					state<=21;
					out<=122;
				end
				if(in == 647) begin
					state<=21;
					out<=123;
				end
				if(in == 648) begin
					state<=21;
					out<=124;
				end
				if(in == 649) begin
					state<=21;
					out<=125;
				end
				if(in == 650) begin
					state<=21;
					out<=126;
				end
				if(in == 651) begin
					state<=21;
					out<=127;
				end
				if(in == 652) begin
					state<=21;
					out<=128;
				end
				if(in == 653) begin
					state<=21;
					out<=129;
				end
				if(in == 654) begin
					state<=21;
					out<=130;
				end
				if(in == 655) begin
					state<=21;
					out<=131;
				end
				if(in == 656) begin
					state<=21;
					out<=132;
				end
				if(in == 657) begin
					state<=21;
					out<=133;
				end
				if(in == 658) begin
					state<=21;
					out<=134;
				end
				if(in == 659) begin
					state<=21;
					out<=135;
				end
				if(in == 660) begin
					state<=21;
					out<=136;
				end
				if(in == 661) begin
					state<=21;
					out<=137;
				end
				if(in == 662) begin
					state<=21;
					out<=138;
				end
				if(in == 663) begin
					state<=21;
					out<=139;
				end
				if(in == 664) begin
					state<=21;
					out<=140;
				end
				if(in == 665) begin
					state<=21;
					out<=141;
				end
				if(in == 666) begin
					state<=21;
					out<=142;
				end
				if(in == 667) begin
					state<=21;
					out<=143;
				end
				if(in == 668) begin
					state<=21;
					out<=144;
				end
				if(in == 669) begin
					state<=21;
					out<=145;
				end
				if(in == 670) begin
					state<=21;
					out<=146;
				end
				if(in == 671) begin
					state<=21;
					out<=147;
				end
				if(in == 672) begin
					state<=21;
					out<=148;
				end
				if(in == 673) begin
					state<=21;
					out<=149;
				end
				if(in == 674) begin
					state<=21;
					out<=150;
				end
				if(in == 675) begin
					state<=21;
					out<=151;
				end
				if(in == 676) begin
					state<=21;
					out<=152;
				end
				if(in == 677) begin
					state<=21;
					out<=153;
				end
				if(in == 678) begin
					state<=21;
					out<=154;
				end
				if(in == 679) begin
					state<=21;
					out<=155;
				end
				if(in == 680) begin
					state<=21;
					out<=156;
				end
				if(in == 681) begin
					state<=21;
					out<=157;
				end
				if(in == 682) begin
					state<=21;
					out<=158;
				end
				if(in == 683) begin
					state<=21;
					out<=159;
				end
				if(in == 684) begin
					state<=21;
					out<=160;
				end
				if(in == 685) begin
					state<=2;
					out<=161;
				end
				if(in == 686) begin
					state<=2;
					out<=162;
				end
				if(in == 687) begin
					state<=2;
					out<=163;
				end
				if(in == 688) begin
					state<=2;
					out<=164;
				end
				if(in == 689) begin
					state<=2;
					out<=165;
				end
				if(in == 690) begin
					state<=2;
					out<=166;
				end
				if(in == 691) begin
					state<=2;
					out<=167;
				end
				if(in == 692) begin
					state<=2;
					out<=168;
				end
				if(in == 693) begin
					state<=2;
					out<=169;
				end
				if(in == 694) begin
					state<=2;
					out<=170;
				end
				if(in == 695) begin
					state<=2;
					out<=171;
				end
				if(in == 696) begin
					state<=2;
					out<=172;
				end
				if(in == 697) begin
					state<=3;
					out<=173;
				end
				if(in == 698) begin
					state<=20;
					out<=174;
				end
				if(in == 699) begin
					state<=3;
					out<=175;
				end
				if(in == 700) begin
					state<=21;
					out<=176;
				end
				if(in == 701) begin
					state<=3;
					out<=177;
				end
				if(in == 702) begin
					state<=21;
					out<=178;
				end
				if(in == 703) begin
					state<=21;
					out<=179;
				end
				if(in == 704) begin
					state<=21;
					out<=180;
				end
				if(in == 705) begin
					state<=21;
					out<=181;
				end
				if(in == 706) begin
					state<=21;
					out<=182;
				end
				if(in == 707) begin
					state<=21;
					out<=183;
				end
				if(in == 708) begin
					state<=21;
					out<=184;
				end
				if(in == 709) begin
					state<=21;
					out<=185;
				end
				if(in == 710) begin
					state<=21;
					out<=186;
				end
				if(in == 711) begin
					state<=21;
					out<=187;
				end
				if(in == 712) begin
					state<=21;
					out<=188;
				end
				if(in == 713) begin
					state<=21;
					out<=189;
				end
				if(in == 714) begin
					state<=21;
					out<=190;
				end
				if(in == 715) begin
					state<=21;
					out<=191;
				end
				if(in == 716) begin
					state<=21;
					out<=192;
				end
				if(in == 717) begin
					state<=21;
					out<=193;
				end
				if(in == 718) begin
					state<=21;
					out<=194;
				end
				if(in == 719) begin
					state<=21;
					out<=195;
				end
				if(in == 720) begin
					state<=21;
					out<=196;
				end
				if(in == 721) begin
					state<=21;
					out<=197;
				end
				if(in == 722) begin
					state<=21;
					out<=198;
				end
				if(in == 723) begin
					state<=21;
					out<=199;
				end
				if(in == 724) begin
					state<=21;
					out<=200;
				end
				if(in == 725) begin
					state<=21;
					out<=201;
				end
				if(in == 726) begin
					state<=21;
					out<=202;
				end
				if(in == 727) begin
					state<=21;
					out<=203;
				end
				if(in == 728) begin
					state<=21;
					out<=204;
				end
				if(in == 729) begin
					state<=21;
					out<=205;
				end
				if(in == 730) begin
					state<=21;
					out<=206;
				end
				if(in == 731) begin
					state<=21;
					out<=207;
				end
				if(in == 732) begin
					state<=21;
					out<=208;
				end
				if(in == 733) begin
					state<=21;
					out<=209;
				end
				if(in == 734) begin
					state<=21;
					out<=210;
				end
				if(in == 735) begin
					state<=21;
					out<=211;
				end
				if(in == 736) begin
					state<=21;
					out<=212;
				end
				if(in == 737) begin
					state<=21;
					out<=213;
				end
				if(in == 738) begin
					state<=21;
					out<=214;
				end
				if(in == 739) begin
					state<=21;
					out<=215;
				end
				if(in == 740) begin
					state<=21;
					out<=216;
				end
				if(in == 741) begin
					state<=21;
					out<=217;
				end
				if(in == 742) begin
					state<=21;
					out<=218;
				end
				if(in == 743) begin
					state<=21;
					out<=219;
				end
				if(in == 744) begin
					state<=21;
					out<=220;
				end
				if(in == 745) begin
					state<=21;
					out<=221;
				end
				if(in == 746) begin
					state<=21;
					out<=222;
				end
				if(in == 747) begin
					state<=21;
					out<=223;
				end
				if(in == 748) begin
					state<=21;
					out<=224;
				end
				if(in == 749) begin
					state<=3;
					out<=225;
				end
				if(in == 750) begin
					state<=20;
					out<=226;
				end
				if(in == 751) begin
					state<=3;
					out<=227;
				end
				if(in == 752) begin
					state<=21;
					out<=228;
				end
				if(in == 753) begin
					state<=3;
					out<=229;
				end
				if(in == 754) begin
					state<=21;
					out<=230;
				end
				if(in == 755) begin
					state<=21;
					out<=231;
				end
				if(in == 756) begin
					state<=21;
					out<=232;
				end
				if(in == 757) begin
					state<=21;
					out<=233;
				end
				if(in == 758) begin
					state<=21;
					out<=234;
				end
				if(in == 759) begin
					state<=21;
					out<=235;
				end
				if(in == 760) begin
					state<=21;
					out<=236;
				end
				if(in == 761) begin
					state<=21;
					out<=237;
				end
				if(in == 762) begin
					state<=21;
					out<=238;
				end
				if(in == 763) begin
					state<=21;
					out<=239;
				end
				if(in == 764) begin
					state<=21;
					out<=240;
				end
				if(in == 765) begin
					state<=21;
					out<=241;
				end
				if(in == 766) begin
					state<=21;
					out<=242;
				end
				if(in == 767) begin
					state<=21;
					out<=243;
				end
				if(in == 768) begin
					state<=21;
					out<=244;
				end
				if(in == 769) begin
					state<=21;
					out<=245;
				end
				if(in == 770) begin
					state<=21;
					out<=246;
				end
				if(in == 771) begin
					state<=21;
					out<=247;
				end
				if(in == 772) begin
					state<=21;
					out<=248;
				end
				if(in == 773) begin
					state<=21;
					out<=249;
				end
				if(in == 774) begin
					state<=21;
					out<=250;
				end
				if(in == 775) begin
					state<=21;
					out<=251;
				end
				if(in == 776) begin
					state<=21;
					out<=252;
				end
				if(in == 777) begin
					state<=21;
					out<=253;
				end
				if(in == 778) begin
					state<=21;
					out<=254;
				end
				if(in == 779) begin
					state<=21;
					out<=255;
				end
				if(in == 780) begin
					state<=21;
					out<=0;
				end
				if(in == 781) begin
					state<=21;
					out<=1;
				end
				if(in == 782) begin
					state<=21;
					out<=2;
				end
				if(in == 783) begin
					state<=21;
					out<=3;
				end
				if(in == 784) begin
					state<=21;
					out<=4;
				end
				if(in == 785) begin
					state<=21;
					out<=5;
				end
				if(in == 786) begin
					state<=21;
					out<=6;
				end
				if(in == 787) begin
					state<=21;
					out<=7;
				end
				if(in == 788) begin
					state<=21;
					out<=8;
				end
				if(in == 789) begin
					state<=21;
					out<=9;
				end
				if(in == 790) begin
					state<=21;
					out<=10;
				end
				if(in == 791) begin
					state<=21;
					out<=11;
				end
				if(in == 792) begin
					state<=21;
					out<=12;
				end
				if(in == 793) begin
					state<=21;
					out<=13;
				end
				if(in == 794) begin
					state<=21;
					out<=14;
				end
				if(in == 795) begin
					state<=21;
					out<=15;
				end
				if(in == 796) begin
					state<=21;
					out<=16;
				end
				if(in == 797) begin
					state<=21;
					out<=17;
				end
				if(in == 798) begin
					state<=21;
					out<=18;
				end
				if(in == 799) begin
					state<=21;
					out<=19;
				end
				if(in == 800) begin
					state<=21;
					out<=20;
				end
				if(in == 801) begin
					state<=2;
					out<=21;
				end
				if(in == 802) begin
					state<=2;
					out<=22;
				end
				if(in == 803) begin
					state<=2;
					out<=23;
				end
				if(in == 804) begin
					state<=2;
					out<=24;
				end
				if(in == 805) begin
					state<=2;
					out<=25;
				end
				if(in == 806) begin
					state<=2;
					out<=26;
				end
				if(in == 807) begin
					state<=2;
					out<=27;
				end
				if(in == 808) begin
					state<=2;
					out<=28;
				end
				if(in == 809) begin
					state<=2;
					out<=29;
				end
				if(in == 810) begin
					state<=2;
					out<=30;
				end
				if(in == 811) begin
					state<=2;
					out<=31;
				end
				if(in == 812) begin
					state<=2;
					out<=32;
				end
				if(in == 813) begin
					state<=3;
					out<=33;
				end
				if(in == 814) begin
					state<=20;
					out<=34;
				end
				if(in == 815) begin
					state<=3;
					out<=35;
				end
				if(in == 816) begin
					state<=21;
					out<=36;
				end
				if(in == 817) begin
					state<=3;
					out<=37;
				end
				if(in == 818) begin
					state<=21;
					out<=38;
				end
				if(in == 819) begin
					state<=21;
					out<=39;
				end
				if(in == 820) begin
					state<=21;
					out<=40;
				end
				if(in == 821) begin
					state<=21;
					out<=41;
				end
				if(in == 822) begin
					state<=21;
					out<=42;
				end
				if(in == 823) begin
					state<=21;
					out<=43;
				end
				if(in == 824) begin
					state<=21;
					out<=44;
				end
				if(in == 825) begin
					state<=21;
					out<=45;
				end
				if(in == 826) begin
					state<=21;
					out<=46;
				end
				if(in == 827) begin
					state<=21;
					out<=47;
				end
				if(in == 828) begin
					state<=21;
					out<=48;
				end
				if(in == 829) begin
					state<=21;
					out<=49;
				end
				if(in == 830) begin
					state<=21;
					out<=50;
				end
				if(in == 831) begin
					state<=21;
					out<=51;
				end
				if(in == 832) begin
					state<=21;
					out<=52;
				end
				if(in == 833) begin
					state<=21;
					out<=53;
				end
				if(in == 834) begin
					state<=21;
					out<=54;
				end
				if(in == 835) begin
					state<=21;
					out<=55;
				end
				if(in == 836) begin
					state<=21;
					out<=56;
				end
				if(in == 837) begin
					state<=21;
					out<=57;
				end
				if(in == 838) begin
					state<=21;
					out<=58;
				end
				if(in == 839) begin
					state<=21;
					out<=59;
				end
				if(in == 840) begin
					state<=21;
					out<=60;
				end
				if(in == 841) begin
					state<=21;
					out<=61;
				end
				if(in == 842) begin
					state<=21;
					out<=62;
				end
				if(in == 843) begin
					state<=21;
					out<=63;
				end
				if(in == 844) begin
					state<=21;
					out<=64;
				end
				if(in == 845) begin
					state<=21;
					out<=65;
				end
				if(in == 846) begin
					state<=21;
					out<=66;
				end
				if(in == 847) begin
					state<=21;
					out<=67;
				end
				if(in == 848) begin
					state<=21;
					out<=68;
				end
				if(in == 849) begin
					state<=21;
					out<=69;
				end
				if(in == 850) begin
					state<=21;
					out<=70;
				end
				if(in == 851) begin
					state<=21;
					out<=71;
				end
				if(in == 852) begin
					state<=21;
					out<=72;
				end
				if(in == 853) begin
					state<=21;
					out<=73;
				end
				if(in == 854) begin
					state<=21;
					out<=74;
				end
				if(in == 855) begin
					state<=21;
					out<=75;
				end
				if(in == 856) begin
					state<=21;
					out<=76;
				end
				if(in == 857) begin
					state<=21;
					out<=77;
				end
				if(in == 858) begin
					state<=21;
					out<=78;
				end
				if(in == 859) begin
					state<=21;
					out<=79;
				end
				if(in == 860) begin
					state<=21;
					out<=80;
				end
				if(in == 861) begin
					state<=21;
					out<=81;
				end
				if(in == 862) begin
					state<=21;
					out<=82;
				end
				if(in == 863) begin
					state<=21;
					out<=83;
				end
				if(in == 864) begin
					state<=21;
					out<=84;
				end
				if(in == 865) begin
					state<=3;
					out<=85;
				end
				if(in == 866) begin
					state<=20;
					out<=86;
				end
				if(in == 867) begin
					state<=3;
					out<=87;
				end
				if(in == 868) begin
					state<=21;
					out<=88;
				end
				if(in == 869) begin
					state<=3;
					out<=89;
				end
				if(in == 870) begin
					state<=21;
					out<=90;
				end
				if(in == 871) begin
					state<=21;
					out<=91;
				end
				if(in == 872) begin
					state<=21;
					out<=92;
				end
				if(in == 873) begin
					state<=21;
					out<=93;
				end
				if(in == 874) begin
					state<=21;
					out<=94;
				end
				if(in == 875) begin
					state<=21;
					out<=95;
				end
				if(in == 876) begin
					state<=21;
					out<=96;
				end
				if(in == 877) begin
					state<=21;
					out<=97;
				end
				if(in == 878) begin
					state<=21;
					out<=98;
				end
				if(in == 879) begin
					state<=21;
					out<=99;
				end
				if(in == 880) begin
					state<=21;
					out<=100;
				end
				if(in == 881) begin
					state<=21;
					out<=101;
				end
				if(in == 882) begin
					state<=21;
					out<=102;
				end
				if(in == 883) begin
					state<=21;
					out<=103;
				end
				if(in == 884) begin
					state<=21;
					out<=104;
				end
				if(in == 885) begin
					state<=21;
					out<=105;
				end
				if(in == 886) begin
					state<=21;
					out<=106;
				end
				if(in == 887) begin
					state<=21;
					out<=107;
				end
				if(in == 888) begin
					state<=21;
					out<=108;
				end
				if(in == 889) begin
					state<=21;
					out<=109;
				end
				if(in == 890) begin
					state<=21;
					out<=110;
				end
				if(in == 891) begin
					state<=21;
					out<=111;
				end
				if(in == 892) begin
					state<=21;
					out<=112;
				end
				if(in == 893) begin
					state<=21;
					out<=113;
				end
				if(in == 894) begin
					state<=21;
					out<=114;
				end
				if(in == 895) begin
					state<=21;
					out<=115;
				end
				if(in == 896) begin
					state<=21;
					out<=116;
				end
				if(in == 897) begin
					state<=21;
					out<=117;
				end
				if(in == 898) begin
					state<=21;
					out<=118;
				end
				if(in == 899) begin
					state<=21;
					out<=119;
				end
				if(in == 900) begin
					state<=21;
					out<=120;
				end
				if(in == 901) begin
					state<=21;
					out<=121;
				end
				if(in == 902) begin
					state<=21;
					out<=122;
				end
				if(in == 903) begin
					state<=21;
					out<=123;
				end
				if(in == 904) begin
					state<=21;
					out<=124;
				end
				if(in == 905) begin
					state<=21;
					out<=125;
				end
				if(in == 906) begin
					state<=21;
					out<=126;
				end
				if(in == 907) begin
					state<=21;
					out<=127;
				end
				if(in == 908) begin
					state<=21;
					out<=128;
				end
				if(in == 909) begin
					state<=21;
					out<=129;
				end
				if(in == 910) begin
					state<=21;
					out<=130;
				end
				if(in == 911) begin
					state<=21;
					out<=131;
				end
				if(in == 912) begin
					state<=21;
					out<=132;
				end
				if(in == 913) begin
					state<=21;
					out<=133;
				end
				if(in == 914) begin
					state<=21;
					out<=134;
				end
				if(in == 915) begin
					state<=21;
					out<=135;
				end
				if(in == 916) begin
					state<=21;
					out<=136;
				end
				if(in == 917) begin
					state<=2;
					out<=137;
				end
				if(in == 918) begin
					state<=2;
					out<=138;
				end
				if(in == 919) begin
					state<=2;
					out<=139;
				end
				if(in == 920) begin
					state<=2;
					out<=140;
				end
				if(in == 921) begin
					state<=2;
					out<=141;
				end
				if(in == 922) begin
					state<=2;
					out<=142;
				end
				if(in == 923) begin
					state<=2;
					out<=143;
				end
				if(in == 924) begin
					state<=2;
					out<=144;
				end
				if(in == 925) begin
					state<=2;
					out<=145;
				end
				if(in == 926) begin
					state<=2;
					out<=146;
				end
				if(in == 927) begin
					state<=2;
					out<=147;
				end
				if(in == 928) begin
					state<=2;
					out<=148;
				end
			end
			21: begin
				if(in == 0) begin
					state<=3;
					out<=149;
				end
				if(in == 1) begin
					state<=1;
					out<=150;
				end
				if(in == 2) begin
					state<=21;
					out<=151;
				end
				if(in == 3) begin
					state<=3;
					out<=152;
				end
				if(in == 4) begin
					state<=22;
					out<=153;
				end
				if(in == 5) begin
					state<=3;
					out<=154;
				end
				if(in == 6) begin
					state<=22;
					out<=155;
				end
				if(in == 7) begin
					state<=22;
					out<=156;
				end
				if(in == 8) begin
					state<=22;
					out<=157;
				end
				if(in == 9) begin
					state<=22;
					out<=158;
				end
				if(in == 10) begin
					state<=22;
					out<=159;
				end
				if(in == 11) begin
					state<=22;
					out<=160;
				end
				if(in == 12) begin
					state<=22;
					out<=161;
				end
				if(in == 13) begin
					state<=22;
					out<=162;
				end
				if(in == 14) begin
					state<=22;
					out<=163;
				end
				if(in == 15) begin
					state<=22;
					out<=164;
				end
				if(in == 16) begin
					state<=22;
					out<=165;
				end
				if(in == 17) begin
					state<=22;
					out<=166;
				end
				if(in == 18) begin
					state<=22;
					out<=167;
				end
				if(in == 19) begin
					state<=22;
					out<=168;
				end
				if(in == 20) begin
					state<=22;
					out<=169;
				end
				if(in == 21) begin
					state<=22;
					out<=170;
				end
				if(in == 22) begin
					state<=22;
					out<=171;
				end
				if(in == 23) begin
					state<=22;
					out<=172;
				end
				if(in == 24) begin
					state<=22;
					out<=173;
				end
				if(in == 25) begin
					state<=22;
					out<=174;
				end
				if(in == 26) begin
					state<=22;
					out<=175;
				end
				if(in == 27) begin
					state<=22;
					out<=176;
				end
				if(in == 28) begin
					state<=22;
					out<=177;
				end
				if(in == 29) begin
					state<=22;
					out<=178;
				end
				if(in == 30) begin
					state<=22;
					out<=179;
				end
				if(in == 31) begin
					state<=22;
					out<=180;
				end
				if(in == 32) begin
					state<=22;
					out<=181;
				end
				if(in == 33) begin
					state<=22;
					out<=182;
				end
				if(in == 34) begin
					state<=22;
					out<=183;
				end
				if(in == 35) begin
					state<=22;
					out<=184;
				end
				if(in == 36) begin
					state<=22;
					out<=185;
				end
				if(in == 37) begin
					state<=22;
					out<=186;
				end
				if(in == 38) begin
					state<=22;
					out<=187;
				end
				if(in == 39) begin
					state<=22;
					out<=188;
				end
				if(in == 40) begin
					state<=22;
					out<=189;
				end
				if(in == 41) begin
					state<=22;
					out<=190;
				end
				if(in == 42) begin
					state<=22;
					out<=191;
				end
				if(in == 43) begin
					state<=22;
					out<=192;
				end
				if(in == 44) begin
					state<=22;
					out<=193;
				end
				if(in == 45) begin
					state<=22;
					out<=194;
				end
				if(in == 46) begin
					state<=22;
					out<=195;
				end
				if(in == 47) begin
					state<=22;
					out<=196;
				end
				if(in == 48) begin
					state<=22;
					out<=197;
				end
				if(in == 49) begin
					state<=22;
					out<=198;
				end
				if(in == 50) begin
					state<=22;
					out<=199;
				end
				if(in == 51) begin
					state<=22;
					out<=200;
				end
				if(in == 52) begin
					state<=22;
					out<=201;
				end
				if(in == 53) begin
					state<=3;
					out<=202;
				end
				if(in == 54) begin
					state<=21;
					out<=203;
				end
				if(in == 55) begin
					state<=3;
					out<=204;
				end
				if(in == 56) begin
					state<=22;
					out<=205;
				end
				if(in == 57) begin
					state<=3;
					out<=206;
				end
				if(in == 58) begin
					state<=22;
					out<=207;
				end
				if(in == 59) begin
					state<=22;
					out<=208;
				end
				if(in == 60) begin
					state<=22;
					out<=209;
				end
				if(in == 61) begin
					state<=22;
					out<=210;
				end
				if(in == 62) begin
					state<=22;
					out<=211;
				end
				if(in == 63) begin
					state<=22;
					out<=212;
				end
				if(in == 64) begin
					state<=22;
					out<=213;
				end
				if(in == 65) begin
					state<=22;
					out<=214;
				end
				if(in == 66) begin
					state<=22;
					out<=215;
				end
				if(in == 67) begin
					state<=22;
					out<=216;
				end
				if(in == 68) begin
					state<=22;
					out<=217;
				end
				if(in == 69) begin
					state<=22;
					out<=218;
				end
				if(in == 70) begin
					state<=22;
					out<=219;
				end
				if(in == 71) begin
					state<=22;
					out<=220;
				end
				if(in == 72) begin
					state<=22;
					out<=221;
				end
				if(in == 73) begin
					state<=22;
					out<=222;
				end
				if(in == 74) begin
					state<=22;
					out<=223;
				end
				if(in == 75) begin
					state<=22;
					out<=224;
				end
				if(in == 76) begin
					state<=22;
					out<=225;
				end
				if(in == 77) begin
					state<=22;
					out<=226;
				end
				if(in == 78) begin
					state<=22;
					out<=227;
				end
				if(in == 79) begin
					state<=22;
					out<=228;
				end
				if(in == 80) begin
					state<=22;
					out<=229;
				end
				if(in == 81) begin
					state<=22;
					out<=230;
				end
				if(in == 82) begin
					state<=22;
					out<=231;
				end
				if(in == 83) begin
					state<=22;
					out<=232;
				end
				if(in == 84) begin
					state<=22;
					out<=233;
				end
				if(in == 85) begin
					state<=22;
					out<=234;
				end
				if(in == 86) begin
					state<=22;
					out<=235;
				end
				if(in == 87) begin
					state<=22;
					out<=236;
				end
				if(in == 88) begin
					state<=22;
					out<=237;
				end
				if(in == 89) begin
					state<=22;
					out<=238;
				end
				if(in == 90) begin
					state<=22;
					out<=239;
				end
				if(in == 91) begin
					state<=22;
					out<=240;
				end
				if(in == 92) begin
					state<=22;
					out<=241;
				end
				if(in == 93) begin
					state<=22;
					out<=242;
				end
				if(in == 94) begin
					state<=22;
					out<=243;
				end
				if(in == 95) begin
					state<=22;
					out<=244;
				end
				if(in == 96) begin
					state<=22;
					out<=245;
				end
				if(in == 97) begin
					state<=22;
					out<=246;
				end
				if(in == 98) begin
					state<=22;
					out<=247;
				end
				if(in == 99) begin
					state<=22;
					out<=248;
				end
				if(in == 100) begin
					state<=22;
					out<=249;
				end
				if(in == 101) begin
					state<=22;
					out<=250;
				end
				if(in == 102) begin
					state<=22;
					out<=251;
				end
				if(in == 103) begin
					state<=22;
					out<=252;
				end
				if(in == 104) begin
					state<=22;
					out<=253;
				end
				if(in == 105) begin
					state<=2;
					out<=254;
				end
				if(in == 106) begin
					state<=2;
					out<=255;
				end
				if(in == 107) begin
					state<=2;
					out<=0;
				end
				if(in == 108) begin
					state<=2;
					out<=1;
				end
				if(in == 109) begin
					state<=2;
					out<=2;
				end
				if(in == 110) begin
					state<=2;
					out<=3;
				end
				if(in == 111) begin
					state<=2;
					out<=4;
				end
				if(in == 112) begin
					state<=2;
					out<=5;
				end
				if(in == 113) begin
					state<=2;
					out<=6;
				end
				if(in == 114) begin
					state<=2;
					out<=7;
				end
				if(in == 115) begin
					state<=2;
					out<=8;
				end
				if(in == 116) begin
					state<=2;
					out<=9;
				end
				if(in == 117) begin
					state<=3;
					out<=10;
				end
				if(in == 118) begin
					state<=21;
					out<=11;
				end
				if(in == 119) begin
					state<=3;
					out<=12;
				end
				if(in == 120) begin
					state<=22;
					out<=13;
				end
				if(in == 121) begin
					state<=3;
					out<=14;
				end
				if(in == 122) begin
					state<=22;
					out<=15;
				end
				if(in == 123) begin
					state<=22;
					out<=16;
				end
				if(in == 124) begin
					state<=22;
					out<=17;
				end
				if(in == 125) begin
					state<=22;
					out<=18;
				end
				if(in == 126) begin
					state<=22;
					out<=19;
				end
				if(in == 127) begin
					state<=22;
					out<=20;
				end
				if(in == 128) begin
					state<=22;
					out<=21;
				end
				if(in == 129) begin
					state<=22;
					out<=22;
				end
				if(in == 130) begin
					state<=22;
					out<=23;
				end
				if(in == 131) begin
					state<=22;
					out<=24;
				end
				if(in == 132) begin
					state<=22;
					out<=25;
				end
				if(in == 133) begin
					state<=22;
					out<=26;
				end
				if(in == 134) begin
					state<=22;
					out<=27;
				end
				if(in == 135) begin
					state<=22;
					out<=28;
				end
				if(in == 136) begin
					state<=22;
					out<=29;
				end
				if(in == 137) begin
					state<=22;
					out<=30;
				end
				if(in == 138) begin
					state<=22;
					out<=31;
				end
				if(in == 139) begin
					state<=22;
					out<=32;
				end
				if(in == 140) begin
					state<=22;
					out<=33;
				end
				if(in == 141) begin
					state<=22;
					out<=34;
				end
				if(in == 142) begin
					state<=22;
					out<=35;
				end
				if(in == 143) begin
					state<=22;
					out<=36;
				end
				if(in == 144) begin
					state<=22;
					out<=37;
				end
				if(in == 145) begin
					state<=22;
					out<=38;
				end
				if(in == 146) begin
					state<=22;
					out<=39;
				end
				if(in == 147) begin
					state<=22;
					out<=40;
				end
				if(in == 148) begin
					state<=22;
					out<=41;
				end
				if(in == 149) begin
					state<=22;
					out<=42;
				end
				if(in == 150) begin
					state<=22;
					out<=43;
				end
				if(in == 151) begin
					state<=22;
					out<=44;
				end
				if(in == 152) begin
					state<=22;
					out<=45;
				end
				if(in == 153) begin
					state<=22;
					out<=46;
				end
				if(in == 154) begin
					state<=22;
					out<=47;
				end
				if(in == 155) begin
					state<=22;
					out<=48;
				end
				if(in == 156) begin
					state<=22;
					out<=49;
				end
				if(in == 157) begin
					state<=22;
					out<=50;
				end
				if(in == 158) begin
					state<=22;
					out<=51;
				end
				if(in == 159) begin
					state<=22;
					out<=52;
				end
				if(in == 160) begin
					state<=22;
					out<=53;
				end
				if(in == 161) begin
					state<=22;
					out<=54;
				end
				if(in == 162) begin
					state<=22;
					out<=55;
				end
				if(in == 163) begin
					state<=22;
					out<=56;
				end
				if(in == 164) begin
					state<=22;
					out<=57;
				end
				if(in == 165) begin
					state<=22;
					out<=58;
				end
				if(in == 166) begin
					state<=22;
					out<=59;
				end
				if(in == 167) begin
					state<=22;
					out<=60;
				end
				if(in == 168) begin
					state<=22;
					out<=61;
				end
				if(in == 169) begin
					state<=3;
					out<=62;
				end
				if(in == 170) begin
					state<=21;
					out<=63;
				end
				if(in == 171) begin
					state<=3;
					out<=64;
				end
				if(in == 172) begin
					state<=22;
					out<=65;
				end
				if(in == 173) begin
					state<=3;
					out<=66;
				end
				if(in == 174) begin
					state<=22;
					out<=67;
				end
				if(in == 175) begin
					state<=22;
					out<=68;
				end
				if(in == 176) begin
					state<=22;
					out<=69;
				end
				if(in == 177) begin
					state<=22;
					out<=70;
				end
				if(in == 178) begin
					state<=22;
					out<=71;
				end
				if(in == 179) begin
					state<=22;
					out<=72;
				end
				if(in == 180) begin
					state<=22;
					out<=73;
				end
				if(in == 181) begin
					state<=22;
					out<=74;
				end
				if(in == 182) begin
					state<=22;
					out<=75;
				end
				if(in == 183) begin
					state<=22;
					out<=76;
				end
				if(in == 184) begin
					state<=22;
					out<=77;
				end
				if(in == 185) begin
					state<=22;
					out<=78;
				end
				if(in == 186) begin
					state<=22;
					out<=79;
				end
				if(in == 187) begin
					state<=22;
					out<=80;
				end
				if(in == 188) begin
					state<=22;
					out<=81;
				end
				if(in == 189) begin
					state<=22;
					out<=82;
				end
				if(in == 190) begin
					state<=22;
					out<=83;
				end
				if(in == 191) begin
					state<=22;
					out<=84;
				end
				if(in == 192) begin
					state<=22;
					out<=85;
				end
				if(in == 193) begin
					state<=22;
					out<=86;
				end
				if(in == 194) begin
					state<=22;
					out<=87;
				end
				if(in == 195) begin
					state<=22;
					out<=88;
				end
				if(in == 196) begin
					state<=22;
					out<=89;
				end
				if(in == 197) begin
					state<=22;
					out<=90;
				end
				if(in == 198) begin
					state<=22;
					out<=91;
				end
				if(in == 199) begin
					state<=22;
					out<=92;
				end
				if(in == 200) begin
					state<=22;
					out<=93;
				end
				if(in == 201) begin
					state<=22;
					out<=94;
				end
				if(in == 202) begin
					state<=22;
					out<=95;
				end
				if(in == 203) begin
					state<=22;
					out<=96;
				end
				if(in == 204) begin
					state<=22;
					out<=97;
				end
				if(in == 205) begin
					state<=22;
					out<=98;
				end
				if(in == 206) begin
					state<=22;
					out<=99;
				end
				if(in == 207) begin
					state<=22;
					out<=100;
				end
				if(in == 208) begin
					state<=22;
					out<=101;
				end
				if(in == 209) begin
					state<=22;
					out<=102;
				end
				if(in == 210) begin
					state<=22;
					out<=103;
				end
				if(in == 211) begin
					state<=22;
					out<=104;
				end
				if(in == 212) begin
					state<=22;
					out<=105;
				end
				if(in == 213) begin
					state<=22;
					out<=106;
				end
				if(in == 214) begin
					state<=22;
					out<=107;
				end
				if(in == 215) begin
					state<=22;
					out<=108;
				end
				if(in == 216) begin
					state<=22;
					out<=109;
				end
				if(in == 217) begin
					state<=22;
					out<=110;
				end
				if(in == 218) begin
					state<=22;
					out<=111;
				end
				if(in == 219) begin
					state<=22;
					out<=112;
				end
				if(in == 220) begin
					state<=22;
					out<=113;
				end
				if(in == 221) begin
					state<=2;
					out<=114;
				end
				if(in == 222) begin
					state<=2;
					out<=115;
				end
				if(in == 223) begin
					state<=2;
					out<=116;
				end
				if(in == 224) begin
					state<=2;
					out<=117;
				end
				if(in == 225) begin
					state<=2;
					out<=118;
				end
				if(in == 226) begin
					state<=2;
					out<=119;
				end
				if(in == 227) begin
					state<=2;
					out<=120;
				end
				if(in == 228) begin
					state<=2;
					out<=121;
				end
				if(in == 229) begin
					state<=2;
					out<=122;
				end
				if(in == 230) begin
					state<=2;
					out<=123;
				end
				if(in == 231) begin
					state<=2;
					out<=124;
				end
				if(in == 232) begin
					state<=2;
					out<=125;
				end
				if(in == 233) begin
					state<=3;
					out<=126;
				end
				if(in == 234) begin
					state<=21;
					out<=127;
				end
				if(in == 235) begin
					state<=3;
					out<=128;
				end
				if(in == 236) begin
					state<=22;
					out<=129;
				end
				if(in == 237) begin
					state<=3;
					out<=130;
				end
				if(in == 238) begin
					state<=22;
					out<=131;
				end
				if(in == 239) begin
					state<=22;
					out<=132;
				end
				if(in == 240) begin
					state<=22;
					out<=133;
				end
				if(in == 241) begin
					state<=22;
					out<=134;
				end
				if(in == 242) begin
					state<=22;
					out<=135;
				end
				if(in == 243) begin
					state<=22;
					out<=136;
				end
				if(in == 244) begin
					state<=22;
					out<=137;
				end
				if(in == 245) begin
					state<=22;
					out<=138;
				end
				if(in == 246) begin
					state<=22;
					out<=139;
				end
				if(in == 247) begin
					state<=22;
					out<=140;
				end
				if(in == 248) begin
					state<=22;
					out<=141;
				end
				if(in == 249) begin
					state<=22;
					out<=142;
				end
				if(in == 250) begin
					state<=22;
					out<=143;
				end
				if(in == 251) begin
					state<=22;
					out<=144;
				end
				if(in == 252) begin
					state<=22;
					out<=145;
				end
				if(in == 253) begin
					state<=22;
					out<=146;
				end
				if(in == 254) begin
					state<=22;
					out<=147;
				end
				if(in == 255) begin
					state<=22;
					out<=148;
				end
				if(in == 256) begin
					state<=22;
					out<=149;
				end
				if(in == 257) begin
					state<=22;
					out<=150;
				end
				if(in == 258) begin
					state<=22;
					out<=151;
				end
				if(in == 259) begin
					state<=22;
					out<=152;
				end
				if(in == 260) begin
					state<=22;
					out<=153;
				end
				if(in == 261) begin
					state<=22;
					out<=154;
				end
				if(in == 262) begin
					state<=22;
					out<=155;
				end
				if(in == 263) begin
					state<=22;
					out<=156;
				end
				if(in == 264) begin
					state<=22;
					out<=157;
				end
				if(in == 265) begin
					state<=22;
					out<=158;
				end
				if(in == 266) begin
					state<=22;
					out<=159;
				end
				if(in == 267) begin
					state<=22;
					out<=160;
				end
				if(in == 268) begin
					state<=22;
					out<=161;
				end
				if(in == 269) begin
					state<=22;
					out<=162;
				end
				if(in == 270) begin
					state<=22;
					out<=163;
				end
				if(in == 271) begin
					state<=22;
					out<=164;
				end
				if(in == 272) begin
					state<=22;
					out<=165;
				end
				if(in == 273) begin
					state<=22;
					out<=166;
				end
				if(in == 274) begin
					state<=22;
					out<=167;
				end
				if(in == 275) begin
					state<=22;
					out<=168;
				end
				if(in == 276) begin
					state<=22;
					out<=169;
				end
				if(in == 277) begin
					state<=22;
					out<=170;
				end
				if(in == 278) begin
					state<=22;
					out<=171;
				end
				if(in == 279) begin
					state<=22;
					out<=172;
				end
				if(in == 280) begin
					state<=22;
					out<=173;
				end
				if(in == 281) begin
					state<=22;
					out<=174;
				end
				if(in == 282) begin
					state<=22;
					out<=175;
				end
				if(in == 283) begin
					state<=22;
					out<=176;
				end
				if(in == 284) begin
					state<=22;
					out<=177;
				end
				if(in == 285) begin
					state<=3;
					out<=178;
				end
				if(in == 286) begin
					state<=21;
					out<=179;
				end
				if(in == 287) begin
					state<=3;
					out<=180;
				end
				if(in == 288) begin
					state<=22;
					out<=181;
				end
				if(in == 289) begin
					state<=3;
					out<=182;
				end
				if(in == 290) begin
					state<=22;
					out<=183;
				end
				if(in == 291) begin
					state<=22;
					out<=184;
				end
				if(in == 292) begin
					state<=22;
					out<=185;
				end
				if(in == 293) begin
					state<=22;
					out<=186;
				end
				if(in == 294) begin
					state<=22;
					out<=187;
				end
				if(in == 295) begin
					state<=22;
					out<=188;
				end
				if(in == 296) begin
					state<=22;
					out<=189;
				end
				if(in == 297) begin
					state<=22;
					out<=190;
				end
				if(in == 298) begin
					state<=22;
					out<=191;
				end
				if(in == 299) begin
					state<=22;
					out<=192;
				end
				if(in == 300) begin
					state<=22;
					out<=193;
				end
				if(in == 301) begin
					state<=22;
					out<=194;
				end
				if(in == 302) begin
					state<=22;
					out<=195;
				end
				if(in == 303) begin
					state<=22;
					out<=196;
				end
				if(in == 304) begin
					state<=22;
					out<=197;
				end
				if(in == 305) begin
					state<=22;
					out<=198;
				end
				if(in == 306) begin
					state<=22;
					out<=199;
				end
				if(in == 307) begin
					state<=22;
					out<=200;
				end
				if(in == 308) begin
					state<=22;
					out<=201;
				end
				if(in == 309) begin
					state<=22;
					out<=202;
				end
				if(in == 310) begin
					state<=22;
					out<=203;
				end
				if(in == 311) begin
					state<=22;
					out<=204;
				end
				if(in == 312) begin
					state<=22;
					out<=205;
				end
				if(in == 313) begin
					state<=22;
					out<=206;
				end
				if(in == 314) begin
					state<=22;
					out<=207;
				end
				if(in == 315) begin
					state<=22;
					out<=208;
				end
				if(in == 316) begin
					state<=22;
					out<=209;
				end
				if(in == 317) begin
					state<=22;
					out<=210;
				end
				if(in == 318) begin
					state<=22;
					out<=211;
				end
				if(in == 319) begin
					state<=22;
					out<=212;
				end
				if(in == 320) begin
					state<=22;
					out<=213;
				end
				if(in == 321) begin
					state<=22;
					out<=214;
				end
				if(in == 322) begin
					state<=22;
					out<=215;
				end
				if(in == 323) begin
					state<=22;
					out<=216;
				end
				if(in == 324) begin
					state<=22;
					out<=217;
				end
				if(in == 325) begin
					state<=22;
					out<=218;
				end
				if(in == 326) begin
					state<=22;
					out<=219;
				end
				if(in == 327) begin
					state<=22;
					out<=220;
				end
				if(in == 328) begin
					state<=22;
					out<=221;
				end
				if(in == 329) begin
					state<=22;
					out<=222;
				end
				if(in == 330) begin
					state<=22;
					out<=223;
				end
				if(in == 331) begin
					state<=22;
					out<=224;
				end
				if(in == 332) begin
					state<=22;
					out<=225;
				end
				if(in == 333) begin
					state<=22;
					out<=226;
				end
				if(in == 334) begin
					state<=22;
					out<=227;
				end
				if(in == 335) begin
					state<=22;
					out<=228;
				end
				if(in == 336) begin
					state<=22;
					out<=229;
				end
				if(in == 337) begin
					state<=2;
					out<=230;
				end
				if(in == 338) begin
					state<=2;
					out<=231;
				end
				if(in == 339) begin
					state<=2;
					out<=232;
				end
				if(in == 340) begin
					state<=2;
					out<=233;
				end
				if(in == 341) begin
					state<=2;
					out<=234;
				end
				if(in == 342) begin
					state<=2;
					out<=235;
				end
				if(in == 343) begin
					state<=2;
					out<=236;
				end
				if(in == 344) begin
					state<=2;
					out<=237;
				end
				if(in == 345) begin
					state<=2;
					out<=238;
				end
				if(in == 346) begin
					state<=2;
					out<=239;
				end
				if(in == 347) begin
					state<=2;
					out<=240;
				end
				if(in == 348) begin
					state<=2;
					out<=241;
				end
				if(in == 349) begin
					state<=3;
					out<=242;
				end
				if(in == 350) begin
					state<=21;
					out<=243;
				end
				if(in == 351) begin
					state<=3;
					out<=244;
				end
				if(in == 352) begin
					state<=22;
					out<=245;
				end
				if(in == 353) begin
					state<=3;
					out<=246;
				end
				if(in == 354) begin
					state<=22;
					out<=247;
				end
				if(in == 355) begin
					state<=22;
					out<=248;
				end
				if(in == 356) begin
					state<=22;
					out<=249;
				end
				if(in == 357) begin
					state<=22;
					out<=250;
				end
				if(in == 358) begin
					state<=22;
					out<=251;
				end
				if(in == 359) begin
					state<=22;
					out<=252;
				end
				if(in == 360) begin
					state<=22;
					out<=253;
				end
				if(in == 361) begin
					state<=22;
					out<=254;
				end
				if(in == 362) begin
					state<=22;
					out<=255;
				end
				if(in == 363) begin
					state<=22;
					out<=0;
				end
				if(in == 364) begin
					state<=22;
					out<=1;
				end
				if(in == 365) begin
					state<=22;
					out<=2;
				end
				if(in == 366) begin
					state<=22;
					out<=3;
				end
				if(in == 367) begin
					state<=22;
					out<=4;
				end
				if(in == 368) begin
					state<=22;
					out<=5;
				end
				if(in == 369) begin
					state<=22;
					out<=6;
				end
				if(in == 370) begin
					state<=22;
					out<=7;
				end
				if(in == 371) begin
					state<=22;
					out<=8;
				end
				if(in == 372) begin
					state<=22;
					out<=9;
				end
				if(in == 373) begin
					state<=22;
					out<=10;
				end
				if(in == 374) begin
					state<=22;
					out<=11;
				end
				if(in == 375) begin
					state<=22;
					out<=12;
				end
				if(in == 376) begin
					state<=22;
					out<=13;
				end
				if(in == 377) begin
					state<=22;
					out<=14;
				end
				if(in == 378) begin
					state<=22;
					out<=15;
				end
				if(in == 379) begin
					state<=22;
					out<=16;
				end
				if(in == 380) begin
					state<=22;
					out<=17;
				end
				if(in == 381) begin
					state<=22;
					out<=18;
				end
				if(in == 382) begin
					state<=22;
					out<=19;
				end
				if(in == 383) begin
					state<=22;
					out<=20;
				end
				if(in == 384) begin
					state<=22;
					out<=21;
				end
				if(in == 385) begin
					state<=22;
					out<=22;
				end
				if(in == 386) begin
					state<=22;
					out<=23;
				end
				if(in == 387) begin
					state<=22;
					out<=24;
				end
				if(in == 388) begin
					state<=22;
					out<=25;
				end
				if(in == 389) begin
					state<=22;
					out<=26;
				end
				if(in == 390) begin
					state<=22;
					out<=27;
				end
				if(in == 391) begin
					state<=22;
					out<=28;
				end
				if(in == 392) begin
					state<=22;
					out<=29;
				end
				if(in == 393) begin
					state<=22;
					out<=30;
				end
				if(in == 394) begin
					state<=22;
					out<=31;
				end
				if(in == 395) begin
					state<=22;
					out<=32;
				end
				if(in == 396) begin
					state<=22;
					out<=33;
				end
				if(in == 397) begin
					state<=22;
					out<=34;
				end
				if(in == 398) begin
					state<=22;
					out<=35;
				end
				if(in == 399) begin
					state<=22;
					out<=36;
				end
				if(in == 400) begin
					state<=22;
					out<=37;
				end
				if(in == 401) begin
					state<=3;
					out<=38;
				end
				if(in == 402) begin
					state<=21;
					out<=39;
				end
				if(in == 403) begin
					state<=3;
					out<=40;
				end
				if(in == 404) begin
					state<=22;
					out<=41;
				end
				if(in == 405) begin
					state<=3;
					out<=42;
				end
				if(in == 406) begin
					state<=22;
					out<=43;
				end
				if(in == 407) begin
					state<=22;
					out<=44;
				end
				if(in == 408) begin
					state<=22;
					out<=45;
				end
				if(in == 409) begin
					state<=22;
					out<=46;
				end
				if(in == 410) begin
					state<=22;
					out<=47;
				end
				if(in == 411) begin
					state<=22;
					out<=48;
				end
				if(in == 412) begin
					state<=22;
					out<=49;
				end
				if(in == 413) begin
					state<=22;
					out<=50;
				end
				if(in == 414) begin
					state<=22;
					out<=51;
				end
				if(in == 415) begin
					state<=22;
					out<=52;
				end
				if(in == 416) begin
					state<=22;
					out<=53;
				end
				if(in == 417) begin
					state<=22;
					out<=54;
				end
				if(in == 418) begin
					state<=22;
					out<=55;
				end
				if(in == 419) begin
					state<=22;
					out<=56;
				end
				if(in == 420) begin
					state<=22;
					out<=57;
				end
				if(in == 421) begin
					state<=22;
					out<=58;
				end
				if(in == 422) begin
					state<=22;
					out<=59;
				end
				if(in == 423) begin
					state<=22;
					out<=60;
				end
				if(in == 424) begin
					state<=22;
					out<=61;
				end
				if(in == 425) begin
					state<=22;
					out<=62;
				end
				if(in == 426) begin
					state<=22;
					out<=63;
				end
				if(in == 427) begin
					state<=22;
					out<=64;
				end
				if(in == 428) begin
					state<=22;
					out<=65;
				end
				if(in == 429) begin
					state<=22;
					out<=66;
				end
				if(in == 430) begin
					state<=22;
					out<=67;
				end
				if(in == 431) begin
					state<=22;
					out<=68;
				end
				if(in == 432) begin
					state<=22;
					out<=69;
				end
				if(in == 433) begin
					state<=22;
					out<=70;
				end
				if(in == 434) begin
					state<=22;
					out<=71;
				end
				if(in == 435) begin
					state<=22;
					out<=72;
				end
				if(in == 436) begin
					state<=22;
					out<=73;
				end
				if(in == 437) begin
					state<=22;
					out<=74;
				end
				if(in == 438) begin
					state<=22;
					out<=75;
				end
				if(in == 439) begin
					state<=22;
					out<=76;
				end
				if(in == 440) begin
					state<=22;
					out<=77;
				end
				if(in == 441) begin
					state<=22;
					out<=78;
				end
				if(in == 442) begin
					state<=22;
					out<=79;
				end
				if(in == 443) begin
					state<=22;
					out<=80;
				end
				if(in == 444) begin
					state<=22;
					out<=81;
				end
				if(in == 445) begin
					state<=22;
					out<=82;
				end
				if(in == 446) begin
					state<=22;
					out<=83;
				end
				if(in == 447) begin
					state<=22;
					out<=84;
				end
				if(in == 448) begin
					state<=22;
					out<=85;
				end
				if(in == 449) begin
					state<=22;
					out<=86;
				end
				if(in == 450) begin
					state<=22;
					out<=87;
				end
				if(in == 451) begin
					state<=22;
					out<=88;
				end
				if(in == 452) begin
					state<=22;
					out<=89;
				end
				if(in == 453) begin
					state<=2;
					out<=90;
				end
				if(in == 454) begin
					state<=2;
					out<=91;
				end
				if(in == 455) begin
					state<=2;
					out<=92;
				end
				if(in == 456) begin
					state<=2;
					out<=93;
				end
				if(in == 457) begin
					state<=2;
					out<=94;
				end
				if(in == 458) begin
					state<=2;
					out<=95;
				end
				if(in == 459) begin
					state<=2;
					out<=96;
				end
				if(in == 460) begin
					state<=2;
					out<=97;
				end
				if(in == 461) begin
					state<=2;
					out<=98;
				end
				if(in == 462) begin
					state<=2;
					out<=99;
				end
				if(in == 463) begin
					state<=2;
					out<=100;
				end
				if(in == 464) begin
					state<=2;
					out<=101;
				end
				if(in == 465) begin
					state<=3;
					out<=102;
				end
				if(in == 466) begin
					state<=21;
					out<=103;
				end
				if(in == 467) begin
					state<=3;
					out<=104;
				end
				if(in == 468) begin
					state<=22;
					out<=105;
				end
				if(in == 469) begin
					state<=3;
					out<=106;
				end
				if(in == 470) begin
					state<=22;
					out<=107;
				end
				if(in == 471) begin
					state<=22;
					out<=108;
				end
				if(in == 472) begin
					state<=22;
					out<=109;
				end
				if(in == 473) begin
					state<=22;
					out<=110;
				end
				if(in == 474) begin
					state<=22;
					out<=111;
				end
				if(in == 475) begin
					state<=22;
					out<=112;
				end
				if(in == 476) begin
					state<=22;
					out<=113;
				end
				if(in == 477) begin
					state<=22;
					out<=114;
				end
				if(in == 478) begin
					state<=22;
					out<=115;
				end
				if(in == 479) begin
					state<=22;
					out<=116;
				end
				if(in == 480) begin
					state<=22;
					out<=117;
				end
				if(in == 481) begin
					state<=22;
					out<=118;
				end
				if(in == 482) begin
					state<=22;
					out<=119;
				end
				if(in == 483) begin
					state<=22;
					out<=120;
				end
				if(in == 484) begin
					state<=22;
					out<=121;
				end
				if(in == 485) begin
					state<=22;
					out<=122;
				end
				if(in == 486) begin
					state<=22;
					out<=123;
				end
				if(in == 487) begin
					state<=22;
					out<=124;
				end
				if(in == 488) begin
					state<=22;
					out<=125;
				end
				if(in == 489) begin
					state<=22;
					out<=126;
				end
				if(in == 490) begin
					state<=22;
					out<=127;
				end
				if(in == 491) begin
					state<=22;
					out<=128;
				end
				if(in == 492) begin
					state<=22;
					out<=129;
				end
				if(in == 493) begin
					state<=22;
					out<=130;
				end
				if(in == 494) begin
					state<=22;
					out<=131;
				end
				if(in == 495) begin
					state<=22;
					out<=132;
				end
				if(in == 496) begin
					state<=22;
					out<=133;
				end
				if(in == 497) begin
					state<=22;
					out<=134;
				end
				if(in == 498) begin
					state<=22;
					out<=135;
				end
				if(in == 499) begin
					state<=22;
					out<=136;
				end
				if(in == 500) begin
					state<=22;
					out<=137;
				end
				if(in == 501) begin
					state<=22;
					out<=138;
				end
				if(in == 502) begin
					state<=22;
					out<=139;
				end
				if(in == 503) begin
					state<=22;
					out<=140;
				end
				if(in == 504) begin
					state<=22;
					out<=141;
				end
				if(in == 505) begin
					state<=22;
					out<=142;
				end
				if(in == 506) begin
					state<=22;
					out<=143;
				end
				if(in == 507) begin
					state<=22;
					out<=144;
				end
				if(in == 508) begin
					state<=22;
					out<=145;
				end
				if(in == 509) begin
					state<=22;
					out<=146;
				end
				if(in == 510) begin
					state<=22;
					out<=147;
				end
				if(in == 511) begin
					state<=22;
					out<=148;
				end
				if(in == 512) begin
					state<=22;
					out<=149;
				end
				if(in == 513) begin
					state<=22;
					out<=150;
				end
				if(in == 514) begin
					state<=22;
					out<=151;
				end
				if(in == 515) begin
					state<=22;
					out<=152;
				end
				if(in == 516) begin
					state<=22;
					out<=153;
				end
				if(in == 517) begin
					state<=3;
					out<=154;
				end
				if(in == 518) begin
					state<=21;
					out<=155;
				end
				if(in == 519) begin
					state<=3;
					out<=156;
				end
				if(in == 520) begin
					state<=22;
					out<=157;
				end
				if(in == 521) begin
					state<=3;
					out<=158;
				end
				if(in == 522) begin
					state<=22;
					out<=159;
				end
				if(in == 523) begin
					state<=22;
					out<=160;
				end
				if(in == 524) begin
					state<=22;
					out<=161;
				end
				if(in == 525) begin
					state<=22;
					out<=162;
				end
				if(in == 526) begin
					state<=22;
					out<=163;
				end
				if(in == 527) begin
					state<=22;
					out<=164;
				end
				if(in == 528) begin
					state<=22;
					out<=165;
				end
				if(in == 529) begin
					state<=22;
					out<=166;
				end
				if(in == 530) begin
					state<=22;
					out<=167;
				end
				if(in == 531) begin
					state<=22;
					out<=168;
				end
				if(in == 532) begin
					state<=22;
					out<=169;
				end
				if(in == 533) begin
					state<=22;
					out<=170;
				end
				if(in == 534) begin
					state<=22;
					out<=171;
				end
				if(in == 535) begin
					state<=22;
					out<=172;
				end
				if(in == 536) begin
					state<=22;
					out<=173;
				end
				if(in == 537) begin
					state<=22;
					out<=174;
				end
				if(in == 538) begin
					state<=22;
					out<=175;
				end
				if(in == 539) begin
					state<=22;
					out<=176;
				end
				if(in == 540) begin
					state<=22;
					out<=177;
				end
				if(in == 541) begin
					state<=22;
					out<=178;
				end
				if(in == 542) begin
					state<=22;
					out<=179;
				end
				if(in == 543) begin
					state<=22;
					out<=180;
				end
				if(in == 544) begin
					state<=22;
					out<=181;
				end
				if(in == 545) begin
					state<=22;
					out<=182;
				end
				if(in == 546) begin
					state<=22;
					out<=183;
				end
				if(in == 547) begin
					state<=22;
					out<=184;
				end
				if(in == 548) begin
					state<=22;
					out<=185;
				end
				if(in == 549) begin
					state<=22;
					out<=186;
				end
				if(in == 550) begin
					state<=22;
					out<=187;
				end
				if(in == 551) begin
					state<=22;
					out<=188;
				end
				if(in == 552) begin
					state<=22;
					out<=189;
				end
				if(in == 553) begin
					state<=22;
					out<=190;
				end
				if(in == 554) begin
					state<=22;
					out<=191;
				end
				if(in == 555) begin
					state<=22;
					out<=192;
				end
				if(in == 556) begin
					state<=22;
					out<=193;
				end
				if(in == 557) begin
					state<=22;
					out<=194;
				end
				if(in == 558) begin
					state<=22;
					out<=195;
				end
				if(in == 559) begin
					state<=22;
					out<=196;
				end
				if(in == 560) begin
					state<=22;
					out<=197;
				end
				if(in == 561) begin
					state<=22;
					out<=198;
				end
				if(in == 562) begin
					state<=22;
					out<=199;
				end
				if(in == 563) begin
					state<=22;
					out<=200;
				end
				if(in == 564) begin
					state<=22;
					out<=201;
				end
				if(in == 565) begin
					state<=22;
					out<=202;
				end
				if(in == 566) begin
					state<=22;
					out<=203;
				end
				if(in == 567) begin
					state<=22;
					out<=204;
				end
				if(in == 568) begin
					state<=22;
					out<=205;
				end
				if(in == 569) begin
					state<=2;
					out<=206;
				end
				if(in == 570) begin
					state<=2;
					out<=207;
				end
				if(in == 571) begin
					state<=2;
					out<=208;
				end
				if(in == 572) begin
					state<=2;
					out<=209;
				end
				if(in == 573) begin
					state<=2;
					out<=210;
				end
				if(in == 574) begin
					state<=2;
					out<=211;
				end
				if(in == 575) begin
					state<=2;
					out<=212;
				end
				if(in == 576) begin
					state<=2;
					out<=213;
				end
				if(in == 577) begin
					state<=2;
					out<=214;
				end
				if(in == 578) begin
					state<=2;
					out<=215;
				end
				if(in == 579) begin
					state<=2;
					out<=216;
				end
				if(in == 580) begin
					state<=2;
					out<=217;
				end
				if(in == 581) begin
					state<=3;
					out<=218;
				end
				if(in == 582) begin
					state<=21;
					out<=219;
				end
				if(in == 583) begin
					state<=3;
					out<=220;
				end
				if(in == 584) begin
					state<=22;
					out<=221;
				end
				if(in == 585) begin
					state<=3;
					out<=222;
				end
				if(in == 586) begin
					state<=22;
					out<=223;
				end
				if(in == 587) begin
					state<=22;
					out<=224;
				end
				if(in == 588) begin
					state<=22;
					out<=225;
				end
				if(in == 589) begin
					state<=22;
					out<=226;
				end
				if(in == 590) begin
					state<=22;
					out<=227;
				end
				if(in == 591) begin
					state<=22;
					out<=228;
				end
				if(in == 592) begin
					state<=22;
					out<=229;
				end
				if(in == 593) begin
					state<=22;
					out<=230;
				end
				if(in == 594) begin
					state<=22;
					out<=231;
				end
				if(in == 595) begin
					state<=22;
					out<=232;
				end
				if(in == 596) begin
					state<=22;
					out<=233;
				end
				if(in == 597) begin
					state<=22;
					out<=234;
				end
				if(in == 598) begin
					state<=22;
					out<=235;
				end
				if(in == 599) begin
					state<=22;
					out<=236;
				end
				if(in == 600) begin
					state<=22;
					out<=237;
				end
				if(in == 601) begin
					state<=22;
					out<=238;
				end
				if(in == 602) begin
					state<=22;
					out<=239;
				end
				if(in == 603) begin
					state<=22;
					out<=240;
				end
				if(in == 604) begin
					state<=22;
					out<=241;
				end
				if(in == 605) begin
					state<=22;
					out<=242;
				end
				if(in == 606) begin
					state<=22;
					out<=243;
				end
				if(in == 607) begin
					state<=22;
					out<=244;
				end
				if(in == 608) begin
					state<=22;
					out<=245;
				end
				if(in == 609) begin
					state<=22;
					out<=246;
				end
				if(in == 610) begin
					state<=22;
					out<=247;
				end
				if(in == 611) begin
					state<=22;
					out<=248;
				end
				if(in == 612) begin
					state<=22;
					out<=249;
				end
				if(in == 613) begin
					state<=22;
					out<=250;
				end
				if(in == 614) begin
					state<=22;
					out<=251;
				end
				if(in == 615) begin
					state<=22;
					out<=252;
				end
				if(in == 616) begin
					state<=22;
					out<=253;
				end
				if(in == 617) begin
					state<=22;
					out<=254;
				end
				if(in == 618) begin
					state<=22;
					out<=255;
				end
				if(in == 619) begin
					state<=22;
					out<=0;
				end
				if(in == 620) begin
					state<=22;
					out<=1;
				end
				if(in == 621) begin
					state<=22;
					out<=2;
				end
				if(in == 622) begin
					state<=22;
					out<=3;
				end
				if(in == 623) begin
					state<=22;
					out<=4;
				end
				if(in == 624) begin
					state<=22;
					out<=5;
				end
				if(in == 625) begin
					state<=22;
					out<=6;
				end
				if(in == 626) begin
					state<=22;
					out<=7;
				end
				if(in == 627) begin
					state<=22;
					out<=8;
				end
				if(in == 628) begin
					state<=22;
					out<=9;
				end
				if(in == 629) begin
					state<=22;
					out<=10;
				end
				if(in == 630) begin
					state<=22;
					out<=11;
				end
				if(in == 631) begin
					state<=22;
					out<=12;
				end
				if(in == 632) begin
					state<=22;
					out<=13;
				end
				if(in == 633) begin
					state<=3;
					out<=14;
				end
				if(in == 634) begin
					state<=21;
					out<=15;
				end
				if(in == 635) begin
					state<=3;
					out<=16;
				end
				if(in == 636) begin
					state<=22;
					out<=17;
				end
				if(in == 637) begin
					state<=3;
					out<=18;
				end
				if(in == 638) begin
					state<=22;
					out<=19;
				end
				if(in == 639) begin
					state<=22;
					out<=20;
				end
				if(in == 640) begin
					state<=22;
					out<=21;
				end
				if(in == 641) begin
					state<=22;
					out<=22;
				end
				if(in == 642) begin
					state<=22;
					out<=23;
				end
				if(in == 643) begin
					state<=22;
					out<=24;
				end
				if(in == 644) begin
					state<=22;
					out<=25;
				end
				if(in == 645) begin
					state<=22;
					out<=26;
				end
				if(in == 646) begin
					state<=22;
					out<=27;
				end
				if(in == 647) begin
					state<=22;
					out<=28;
				end
				if(in == 648) begin
					state<=22;
					out<=29;
				end
				if(in == 649) begin
					state<=22;
					out<=30;
				end
				if(in == 650) begin
					state<=22;
					out<=31;
				end
				if(in == 651) begin
					state<=22;
					out<=32;
				end
				if(in == 652) begin
					state<=22;
					out<=33;
				end
				if(in == 653) begin
					state<=22;
					out<=34;
				end
				if(in == 654) begin
					state<=22;
					out<=35;
				end
				if(in == 655) begin
					state<=22;
					out<=36;
				end
				if(in == 656) begin
					state<=22;
					out<=37;
				end
				if(in == 657) begin
					state<=22;
					out<=38;
				end
				if(in == 658) begin
					state<=22;
					out<=39;
				end
				if(in == 659) begin
					state<=22;
					out<=40;
				end
				if(in == 660) begin
					state<=22;
					out<=41;
				end
				if(in == 661) begin
					state<=22;
					out<=42;
				end
				if(in == 662) begin
					state<=22;
					out<=43;
				end
				if(in == 663) begin
					state<=22;
					out<=44;
				end
				if(in == 664) begin
					state<=22;
					out<=45;
				end
				if(in == 665) begin
					state<=22;
					out<=46;
				end
				if(in == 666) begin
					state<=22;
					out<=47;
				end
				if(in == 667) begin
					state<=22;
					out<=48;
				end
				if(in == 668) begin
					state<=22;
					out<=49;
				end
				if(in == 669) begin
					state<=22;
					out<=50;
				end
				if(in == 670) begin
					state<=22;
					out<=51;
				end
				if(in == 671) begin
					state<=22;
					out<=52;
				end
				if(in == 672) begin
					state<=22;
					out<=53;
				end
				if(in == 673) begin
					state<=22;
					out<=54;
				end
				if(in == 674) begin
					state<=22;
					out<=55;
				end
				if(in == 675) begin
					state<=22;
					out<=56;
				end
				if(in == 676) begin
					state<=22;
					out<=57;
				end
				if(in == 677) begin
					state<=22;
					out<=58;
				end
				if(in == 678) begin
					state<=22;
					out<=59;
				end
				if(in == 679) begin
					state<=22;
					out<=60;
				end
				if(in == 680) begin
					state<=22;
					out<=61;
				end
				if(in == 681) begin
					state<=22;
					out<=62;
				end
				if(in == 682) begin
					state<=22;
					out<=63;
				end
				if(in == 683) begin
					state<=22;
					out<=64;
				end
				if(in == 684) begin
					state<=22;
					out<=65;
				end
				if(in == 685) begin
					state<=2;
					out<=66;
				end
				if(in == 686) begin
					state<=2;
					out<=67;
				end
				if(in == 687) begin
					state<=2;
					out<=68;
				end
				if(in == 688) begin
					state<=2;
					out<=69;
				end
				if(in == 689) begin
					state<=2;
					out<=70;
				end
				if(in == 690) begin
					state<=2;
					out<=71;
				end
				if(in == 691) begin
					state<=2;
					out<=72;
				end
				if(in == 692) begin
					state<=2;
					out<=73;
				end
				if(in == 693) begin
					state<=2;
					out<=74;
				end
				if(in == 694) begin
					state<=2;
					out<=75;
				end
				if(in == 695) begin
					state<=2;
					out<=76;
				end
				if(in == 696) begin
					state<=2;
					out<=77;
				end
				if(in == 697) begin
					state<=3;
					out<=78;
				end
				if(in == 698) begin
					state<=21;
					out<=79;
				end
				if(in == 699) begin
					state<=3;
					out<=80;
				end
				if(in == 700) begin
					state<=22;
					out<=81;
				end
				if(in == 701) begin
					state<=3;
					out<=82;
				end
				if(in == 702) begin
					state<=22;
					out<=83;
				end
				if(in == 703) begin
					state<=22;
					out<=84;
				end
				if(in == 704) begin
					state<=22;
					out<=85;
				end
				if(in == 705) begin
					state<=22;
					out<=86;
				end
				if(in == 706) begin
					state<=22;
					out<=87;
				end
				if(in == 707) begin
					state<=22;
					out<=88;
				end
				if(in == 708) begin
					state<=22;
					out<=89;
				end
				if(in == 709) begin
					state<=22;
					out<=90;
				end
				if(in == 710) begin
					state<=22;
					out<=91;
				end
				if(in == 711) begin
					state<=22;
					out<=92;
				end
				if(in == 712) begin
					state<=22;
					out<=93;
				end
				if(in == 713) begin
					state<=22;
					out<=94;
				end
				if(in == 714) begin
					state<=22;
					out<=95;
				end
				if(in == 715) begin
					state<=22;
					out<=96;
				end
				if(in == 716) begin
					state<=22;
					out<=97;
				end
				if(in == 717) begin
					state<=22;
					out<=98;
				end
				if(in == 718) begin
					state<=22;
					out<=99;
				end
				if(in == 719) begin
					state<=22;
					out<=100;
				end
				if(in == 720) begin
					state<=22;
					out<=101;
				end
				if(in == 721) begin
					state<=22;
					out<=102;
				end
				if(in == 722) begin
					state<=22;
					out<=103;
				end
				if(in == 723) begin
					state<=22;
					out<=104;
				end
				if(in == 724) begin
					state<=22;
					out<=105;
				end
				if(in == 725) begin
					state<=22;
					out<=106;
				end
				if(in == 726) begin
					state<=22;
					out<=107;
				end
				if(in == 727) begin
					state<=22;
					out<=108;
				end
				if(in == 728) begin
					state<=22;
					out<=109;
				end
				if(in == 729) begin
					state<=22;
					out<=110;
				end
				if(in == 730) begin
					state<=22;
					out<=111;
				end
				if(in == 731) begin
					state<=22;
					out<=112;
				end
				if(in == 732) begin
					state<=22;
					out<=113;
				end
				if(in == 733) begin
					state<=22;
					out<=114;
				end
				if(in == 734) begin
					state<=22;
					out<=115;
				end
				if(in == 735) begin
					state<=22;
					out<=116;
				end
				if(in == 736) begin
					state<=22;
					out<=117;
				end
				if(in == 737) begin
					state<=22;
					out<=118;
				end
				if(in == 738) begin
					state<=22;
					out<=119;
				end
				if(in == 739) begin
					state<=22;
					out<=120;
				end
				if(in == 740) begin
					state<=22;
					out<=121;
				end
				if(in == 741) begin
					state<=22;
					out<=122;
				end
				if(in == 742) begin
					state<=22;
					out<=123;
				end
				if(in == 743) begin
					state<=22;
					out<=124;
				end
				if(in == 744) begin
					state<=22;
					out<=125;
				end
				if(in == 745) begin
					state<=22;
					out<=126;
				end
				if(in == 746) begin
					state<=22;
					out<=127;
				end
				if(in == 747) begin
					state<=22;
					out<=128;
				end
				if(in == 748) begin
					state<=22;
					out<=129;
				end
				if(in == 749) begin
					state<=3;
					out<=130;
				end
				if(in == 750) begin
					state<=21;
					out<=131;
				end
				if(in == 751) begin
					state<=3;
					out<=132;
				end
				if(in == 752) begin
					state<=22;
					out<=133;
				end
				if(in == 753) begin
					state<=3;
					out<=134;
				end
				if(in == 754) begin
					state<=22;
					out<=135;
				end
				if(in == 755) begin
					state<=22;
					out<=136;
				end
				if(in == 756) begin
					state<=22;
					out<=137;
				end
				if(in == 757) begin
					state<=22;
					out<=138;
				end
				if(in == 758) begin
					state<=22;
					out<=139;
				end
				if(in == 759) begin
					state<=22;
					out<=140;
				end
				if(in == 760) begin
					state<=22;
					out<=141;
				end
				if(in == 761) begin
					state<=22;
					out<=142;
				end
				if(in == 762) begin
					state<=22;
					out<=143;
				end
				if(in == 763) begin
					state<=22;
					out<=144;
				end
				if(in == 764) begin
					state<=22;
					out<=145;
				end
				if(in == 765) begin
					state<=22;
					out<=146;
				end
				if(in == 766) begin
					state<=22;
					out<=147;
				end
				if(in == 767) begin
					state<=22;
					out<=148;
				end
				if(in == 768) begin
					state<=22;
					out<=149;
				end
				if(in == 769) begin
					state<=22;
					out<=150;
				end
				if(in == 770) begin
					state<=22;
					out<=151;
				end
				if(in == 771) begin
					state<=22;
					out<=152;
				end
				if(in == 772) begin
					state<=22;
					out<=153;
				end
				if(in == 773) begin
					state<=22;
					out<=154;
				end
				if(in == 774) begin
					state<=22;
					out<=155;
				end
				if(in == 775) begin
					state<=22;
					out<=156;
				end
				if(in == 776) begin
					state<=22;
					out<=157;
				end
				if(in == 777) begin
					state<=22;
					out<=158;
				end
				if(in == 778) begin
					state<=22;
					out<=159;
				end
				if(in == 779) begin
					state<=22;
					out<=160;
				end
				if(in == 780) begin
					state<=22;
					out<=161;
				end
				if(in == 781) begin
					state<=22;
					out<=162;
				end
				if(in == 782) begin
					state<=22;
					out<=163;
				end
				if(in == 783) begin
					state<=22;
					out<=164;
				end
				if(in == 784) begin
					state<=22;
					out<=165;
				end
				if(in == 785) begin
					state<=22;
					out<=166;
				end
				if(in == 786) begin
					state<=22;
					out<=167;
				end
				if(in == 787) begin
					state<=22;
					out<=168;
				end
				if(in == 788) begin
					state<=22;
					out<=169;
				end
				if(in == 789) begin
					state<=22;
					out<=170;
				end
				if(in == 790) begin
					state<=22;
					out<=171;
				end
				if(in == 791) begin
					state<=22;
					out<=172;
				end
				if(in == 792) begin
					state<=22;
					out<=173;
				end
				if(in == 793) begin
					state<=22;
					out<=174;
				end
				if(in == 794) begin
					state<=22;
					out<=175;
				end
				if(in == 795) begin
					state<=22;
					out<=176;
				end
				if(in == 796) begin
					state<=22;
					out<=177;
				end
				if(in == 797) begin
					state<=22;
					out<=178;
				end
				if(in == 798) begin
					state<=22;
					out<=179;
				end
				if(in == 799) begin
					state<=22;
					out<=180;
				end
				if(in == 800) begin
					state<=22;
					out<=181;
				end
				if(in == 801) begin
					state<=2;
					out<=182;
				end
				if(in == 802) begin
					state<=2;
					out<=183;
				end
				if(in == 803) begin
					state<=2;
					out<=184;
				end
				if(in == 804) begin
					state<=2;
					out<=185;
				end
				if(in == 805) begin
					state<=2;
					out<=186;
				end
				if(in == 806) begin
					state<=2;
					out<=187;
				end
				if(in == 807) begin
					state<=2;
					out<=188;
				end
				if(in == 808) begin
					state<=2;
					out<=189;
				end
				if(in == 809) begin
					state<=2;
					out<=190;
				end
				if(in == 810) begin
					state<=2;
					out<=191;
				end
				if(in == 811) begin
					state<=2;
					out<=192;
				end
				if(in == 812) begin
					state<=2;
					out<=193;
				end
				if(in == 813) begin
					state<=3;
					out<=194;
				end
				if(in == 814) begin
					state<=21;
					out<=195;
				end
				if(in == 815) begin
					state<=3;
					out<=196;
				end
				if(in == 816) begin
					state<=22;
					out<=197;
				end
				if(in == 817) begin
					state<=3;
					out<=198;
				end
				if(in == 818) begin
					state<=22;
					out<=199;
				end
				if(in == 819) begin
					state<=22;
					out<=200;
				end
				if(in == 820) begin
					state<=22;
					out<=201;
				end
				if(in == 821) begin
					state<=22;
					out<=202;
				end
				if(in == 822) begin
					state<=22;
					out<=203;
				end
				if(in == 823) begin
					state<=22;
					out<=204;
				end
				if(in == 824) begin
					state<=22;
					out<=205;
				end
				if(in == 825) begin
					state<=22;
					out<=206;
				end
				if(in == 826) begin
					state<=22;
					out<=207;
				end
				if(in == 827) begin
					state<=22;
					out<=208;
				end
				if(in == 828) begin
					state<=22;
					out<=209;
				end
				if(in == 829) begin
					state<=22;
					out<=210;
				end
				if(in == 830) begin
					state<=22;
					out<=211;
				end
				if(in == 831) begin
					state<=22;
					out<=212;
				end
				if(in == 832) begin
					state<=22;
					out<=213;
				end
				if(in == 833) begin
					state<=22;
					out<=214;
				end
				if(in == 834) begin
					state<=22;
					out<=215;
				end
				if(in == 835) begin
					state<=22;
					out<=216;
				end
				if(in == 836) begin
					state<=22;
					out<=217;
				end
				if(in == 837) begin
					state<=22;
					out<=218;
				end
				if(in == 838) begin
					state<=22;
					out<=219;
				end
				if(in == 839) begin
					state<=22;
					out<=220;
				end
				if(in == 840) begin
					state<=22;
					out<=221;
				end
				if(in == 841) begin
					state<=22;
					out<=222;
				end
				if(in == 842) begin
					state<=22;
					out<=223;
				end
				if(in == 843) begin
					state<=22;
					out<=224;
				end
				if(in == 844) begin
					state<=22;
					out<=225;
				end
				if(in == 845) begin
					state<=22;
					out<=226;
				end
				if(in == 846) begin
					state<=22;
					out<=227;
				end
				if(in == 847) begin
					state<=22;
					out<=228;
				end
				if(in == 848) begin
					state<=22;
					out<=229;
				end
				if(in == 849) begin
					state<=22;
					out<=230;
				end
				if(in == 850) begin
					state<=22;
					out<=231;
				end
				if(in == 851) begin
					state<=22;
					out<=232;
				end
				if(in == 852) begin
					state<=22;
					out<=233;
				end
				if(in == 853) begin
					state<=22;
					out<=234;
				end
				if(in == 854) begin
					state<=22;
					out<=235;
				end
				if(in == 855) begin
					state<=22;
					out<=236;
				end
				if(in == 856) begin
					state<=22;
					out<=237;
				end
				if(in == 857) begin
					state<=22;
					out<=238;
				end
				if(in == 858) begin
					state<=22;
					out<=239;
				end
				if(in == 859) begin
					state<=22;
					out<=240;
				end
				if(in == 860) begin
					state<=22;
					out<=241;
				end
				if(in == 861) begin
					state<=22;
					out<=242;
				end
				if(in == 862) begin
					state<=22;
					out<=243;
				end
				if(in == 863) begin
					state<=22;
					out<=244;
				end
				if(in == 864) begin
					state<=22;
					out<=245;
				end
				if(in == 865) begin
					state<=3;
					out<=246;
				end
				if(in == 866) begin
					state<=21;
					out<=247;
				end
				if(in == 867) begin
					state<=3;
					out<=248;
				end
				if(in == 868) begin
					state<=22;
					out<=249;
				end
				if(in == 869) begin
					state<=3;
					out<=250;
				end
				if(in == 870) begin
					state<=22;
					out<=251;
				end
				if(in == 871) begin
					state<=22;
					out<=252;
				end
				if(in == 872) begin
					state<=22;
					out<=253;
				end
				if(in == 873) begin
					state<=22;
					out<=254;
				end
				if(in == 874) begin
					state<=22;
					out<=255;
				end
				if(in == 875) begin
					state<=22;
					out<=0;
				end
				if(in == 876) begin
					state<=22;
					out<=1;
				end
				if(in == 877) begin
					state<=22;
					out<=2;
				end
				if(in == 878) begin
					state<=22;
					out<=3;
				end
				if(in == 879) begin
					state<=22;
					out<=4;
				end
				if(in == 880) begin
					state<=22;
					out<=5;
				end
				if(in == 881) begin
					state<=22;
					out<=6;
				end
				if(in == 882) begin
					state<=22;
					out<=7;
				end
				if(in == 883) begin
					state<=22;
					out<=8;
				end
				if(in == 884) begin
					state<=22;
					out<=9;
				end
				if(in == 885) begin
					state<=22;
					out<=10;
				end
				if(in == 886) begin
					state<=22;
					out<=11;
				end
				if(in == 887) begin
					state<=22;
					out<=12;
				end
				if(in == 888) begin
					state<=22;
					out<=13;
				end
				if(in == 889) begin
					state<=22;
					out<=14;
				end
				if(in == 890) begin
					state<=22;
					out<=15;
				end
				if(in == 891) begin
					state<=22;
					out<=16;
				end
				if(in == 892) begin
					state<=22;
					out<=17;
				end
				if(in == 893) begin
					state<=22;
					out<=18;
				end
				if(in == 894) begin
					state<=22;
					out<=19;
				end
				if(in == 895) begin
					state<=22;
					out<=20;
				end
				if(in == 896) begin
					state<=22;
					out<=21;
				end
				if(in == 897) begin
					state<=22;
					out<=22;
				end
				if(in == 898) begin
					state<=22;
					out<=23;
				end
				if(in == 899) begin
					state<=22;
					out<=24;
				end
				if(in == 900) begin
					state<=22;
					out<=25;
				end
				if(in == 901) begin
					state<=22;
					out<=26;
				end
				if(in == 902) begin
					state<=22;
					out<=27;
				end
				if(in == 903) begin
					state<=22;
					out<=28;
				end
				if(in == 904) begin
					state<=22;
					out<=29;
				end
				if(in == 905) begin
					state<=22;
					out<=30;
				end
				if(in == 906) begin
					state<=22;
					out<=31;
				end
				if(in == 907) begin
					state<=22;
					out<=32;
				end
				if(in == 908) begin
					state<=22;
					out<=33;
				end
				if(in == 909) begin
					state<=22;
					out<=34;
				end
				if(in == 910) begin
					state<=22;
					out<=35;
				end
				if(in == 911) begin
					state<=22;
					out<=36;
				end
				if(in == 912) begin
					state<=22;
					out<=37;
				end
				if(in == 913) begin
					state<=22;
					out<=38;
				end
				if(in == 914) begin
					state<=22;
					out<=39;
				end
				if(in == 915) begin
					state<=22;
					out<=40;
				end
				if(in == 916) begin
					state<=22;
					out<=41;
				end
				if(in == 917) begin
					state<=2;
					out<=42;
				end
				if(in == 918) begin
					state<=2;
					out<=43;
				end
				if(in == 919) begin
					state<=2;
					out<=44;
				end
				if(in == 920) begin
					state<=2;
					out<=45;
				end
				if(in == 921) begin
					state<=2;
					out<=46;
				end
				if(in == 922) begin
					state<=2;
					out<=47;
				end
				if(in == 923) begin
					state<=2;
					out<=48;
				end
				if(in == 924) begin
					state<=2;
					out<=49;
				end
				if(in == 925) begin
					state<=2;
					out<=50;
				end
				if(in == 926) begin
					state<=2;
					out<=51;
				end
				if(in == 927) begin
					state<=2;
					out<=52;
				end
				if(in == 928) begin
					state<=2;
					out<=53;
				end
			end
			22: begin
				if(in == 0) begin
					state<=13;
					out<=54;
				end
				if(in == 1) begin
					state<=1;
					out<=55;
				end
				if(in == 2) begin
					state<=22;
					out<=56;
				end
				if(in == 3) begin
					state<=13;
					out<=57;
				end
				if(in == 4) begin
					state<=22;
					out<=58;
				end
				if(in == 5) begin
					state<=13;
					out<=59;
				end
				if(in == 6) begin
					state<=22;
					out<=60;
				end
				if(in == 7) begin
					state<=22;
					out<=61;
				end
				if(in == 8) begin
					state<=22;
					out<=62;
				end
				if(in == 9) begin
					state<=22;
					out<=63;
				end
				if(in == 10) begin
					state<=22;
					out<=64;
				end
				if(in == 11) begin
					state<=22;
					out<=65;
				end
				if(in == 12) begin
					state<=22;
					out<=66;
				end
				if(in == 13) begin
					state<=22;
					out<=67;
				end
				if(in == 14) begin
					state<=22;
					out<=68;
				end
				if(in == 15) begin
					state<=22;
					out<=69;
				end
				if(in == 16) begin
					state<=22;
					out<=70;
				end
				if(in == 17) begin
					state<=22;
					out<=71;
				end
				if(in == 18) begin
					state<=22;
					out<=72;
				end
				if(in == 19) begin
					state<=22;
					out<=73;
				end
				if(in == 20) begin
					state<=22;
					out<=74;
				end
				if(in == 21) begin
					state<=22;
					out<=75;
				end
				if(in == 22) begin
					state<=22;
					out<=76;
				end
				if(in == 23) begin
					state<=22;
					out<=77;
				end
				if(in == 24) begin
					state<=22;
					out<=78;
				end
				if(in == 25) begin
					state<=22;
					out<=79;
				end
				if(in == 26) begin
					state<=22;
					out<=80;
				end
				if(in == 27) begin
					state<=22;
					out<=81;
				end
				if(in == 28) begin
					state<=22;
					out<=82;
				end
				if(in == 29) begin
					state<=22;
					out<=83;
				end
				if(in == 30) begin
					state<=22;
					out<=84;
				end
				if(in == 31) begin
					state<=22;
					out<=85;
				end
				if(in == 32) begin
					state<=22;
					out<=86;
				end
				if(in == 33) begin
					state<=22;
					out<=87;
				end
				if(in == 34) begin
					state<=22;
					out<=88;
				end
				if(in == 35) begin
					state<=22;
					out<=89;
				end
				if(in == 36) begin
					state<=22;
					out<=90;
				end
				if(in == 37) begin
					state<=23;
					out<=91;
				end
				if(in == 38) begin
					state<=23;
					out<=92;
				end
				if(in == 39) begin
					state<=23;
					out<=93;
				end
				if(in == 40) begin
					state<=23;
					out<=94;
				end
				if(in == 41) begin
					state<=23;
					out<=95;
				end
				if(in == 42) begin
					state<=23;
					out<=96;
				end
				if(in == 43) begin
					state<=23;
					out<=97;
				end
				if(in == 44) begin
					state<=23;
					out<=98;
				end
				if(in == 45) begin
					state<=23;
					out<=99;
				end
				if(in == 46) begin
					state<=23;
					out<=100;
				end
				if(in == 47) begin
					state<=23;
					out<=101;
				end
				if(in == 48) begin
					state<=23;
					out<=102;
				end
				if(in == 49) begin
					state<=23;
					out<=103;
				end
				if(in == 50) begin
					state<=23;
					out<=104;
				end
				if(in == 51) begin
					state<=23;
					out<=105;
				end
				if(in == 52) begin
					state<=23;
					out<=106;
				end
				if(in == 53) begin
					state<=13;
					out<=107;
				end
				if(in == 54) begin
					state<=22;
					out<=108;
				end
				if(in == 55) begin
					state<=13;
					out<=109;
				end
				if(in == 56) begin
					state<=22;
					out<=110;
				end
				if(in == 57) begin
					state<=13;
					out<=111;
				end
				if(in == 58) begin
					state<=22;
					out<=112;
				end
				if(in == 59) begin
					state<=22;
					out<=113;
				end
				if(in == 60) begin
					state<=22;
					out<=114;
				end
				if(in == 61) begin
					state<=22;
					out<=115;
				end
				if(in == 62) begin
					state<=22;
					out<=116;
				end
				if(in == 63) begin
					state<=22;
					out<=117;
				end
				if(in == 64) begin
					state<=22;
					out<=118;
				end
				if(in == 65) begin
					state<=22;
					out<=119;
				end
				if(in == 66) begin
					state<=22;
					out<=120;
				end
				if(in == 67) begin
					state<=22;
					out<=121;
				end
				if(in == 68) begin
					state<=22;
					out<=122;
				end
				if(in == 69) begin
					state<=22;
					out<=123;
				end
				if(in == 70) begin
					state<=22;
					out<=124;
				end
				if(in == 71) begin
					state<=22;
					out<=125;
				end
				if(in == 72) begin
					state<=22;
					out<=126;
				end
				if(in == 73) begin
					state<=22;
					out<=127;
				end
				if(in == 74) begin
					state<=22;
					out<=128;
				end
				if(in == 75) begin
					state<=22;
					out<=129;
				end
				if(in == 76) begin
					state<=22;
					out<=130;
				end
				if(in == 77) begin
					state<=22;
					out<=131;
				end
				if(in == 78) begin
					state<=22;
					out<=132;
				end
				if(in == 79) begin
					state<=22;
					out<=133;
				end
				if(in == 80) begin
					state<=22;
					out<=134;
				end
				if(in == 81) begin
					state<=22;
					out<=135;
				end
				if(in == 82) begin
					state<=22;
					out<=136;
				end
				if(in == 83) begin
					state<=22;
					out<=137;
				end
				if(in == 84) begin
					state<=22;
					out<=138;
				end
				if(in == 85) begin
					state<=22;
					out<=139;
				end
				if(in == 86) begin
					state<=22;
					out<=140;
				end
				if(in == 87) begin
					state<=22;
					out<=141;
				end
				if(in == 88) begin
					state<=22;
					out<=142;
				end
				if(in == 89) begin
					state<=23;
					out<=143;
				end
				if(in == 90) begin
					state<=23;
					out<=144;
				end
				if(in == 91) begin
					state<=23;
					out<=145;
				end
				if(in == 92) begin
					state<=23;
					out<=146;
				end
				if(in == 93) begin
					state<=23;
					out<=147;
				end
				if(in == 94) begin
					state<=23;
					out<=148;
				end
				if(in == 95) begin
					state<=23;
					out<=149;
				end
				if(in == 96) begin
					state<=23;
					out<=150;
				end
				if(in == 97) begin
					state<=23;
					out<=151;
				end
				if(in == 98) begin
					state<=23;
					out<=152;
				end
				if(in == 99) begin
					state<=23;
					out<=153;
				end
				if(in == 100) begin
					state<=23;
					out<=154;
				end
				if(in == 101) begin
					state<=23;
					out<=155;
				end
				if(in == 102) begin
					state<=23;
					out<=156;
				end
				if(in == 103) begin
					state<=23;
					out<=157;
				end
				if(in == 104) begin
					state<=23;
					out<=158;
				end
				if(in == 105) begin
					state<=2;
					out<=159;
				end
				if(in == 106) begin
					state<=2;
					out<=160;
				end
				if(in == 107) begin
					state<=2;
					out<=161;
				end
				if(in == 108) begin
					state<=2;
					out<=162;
				end
				if(in == 109) begin
					state<=2;
					out<=163;
				end
				if(in == 110) begin
					state<=2;
					out<=164;
				end
				if(in == 111) begin
					state<=2;
					out<=165;
				end
				if(in == 112) begin
					state<=2;
					out<=166;
				end
				if(in == 113) begin
					state<=2;
					out<=167;
				end
				if(in == 114) begin
					state<=2;
					out<=168;
				end
				if(in == 115) begin
					state<=2;
					out<=169;
				end
				if(in == 116) begin
					state<=2;
					out<=170;
				end
				if(in == 117) begin
					state<=13;
					out<=171;
				end
				if(in == 118) begin
					state<=22;
					out<=172;
				end
				if(in == 119) begin
					state<=13;
					out<=173;
				end
				if(in == 120) begin
					state<=22;
					out<=174;
				end
				if(in == 121) begin
					state<=13;
					out<=175;
				end
				if(in == 122) begin
					state<=22;
					out<=176;
				end
				if(in == 123) begin
					state<=22;
					out<=177;
				end
				if(in == 124) begin
					state<=22;
					out<=178;
				end
				if(in == 125) begin
					state<=22;
					out<=179;
				end
				if(in == 126) begin
					state<=22;
					out<=180;
				end
				if(in == 127) begin
					state<=22;
					out<=181;
				end
				if(in == 128) begin
					state<=22;
					out<=182;
				end
				if(in == 129) begin
					state<=22;
					out<=183;
				end
				if(in == 130) begin
					state<=22;
					out<=184;
				end
				if(in == 131) begin
					state<=22;
					out<=185;
				end
				if(in == 132) begin
					state<=22;
					out<=186;
				end
				if(in == 133) begin
					state<=22;
					out<=187;
				end
				if(in == 134) begin
					state<=22;
					out<=188;
				end
				if(in == 135) begin
					state<=22;
					out<=189;
				end
				if(in == 136) begin
					state<=22;
					out<=190;
				end
				if(in == 137) begin
					state<=22;
					out<=191;
				end
				if(in == 138) begin
					state<=22;
					out<=192;
				end
				if(in == 139) begin
					state<=22;
					out<=193;
				end
				if(in == 140) begin
					state<=22;
					out<=194;
				end
				if(in == 141) begin
					state<=22;
					out<=195;
				end
				if(in == 142) begin
					state<=22;
					out<=196;
				end
				if(in == 143) begin
					state<=22;
					out<=197;
				end
				if(in == 144) begin
					state<=22;
					out<=198;
				end
				if(in == 145) begin
					state<=22;
					out<=199;
				end
				if(in == 146) begin
					state<=22;
					out<=200;
				end
				if(in == 147) begin
					state<=22;
					out<=201;
				end
				if(in == 148) begin
					state<=22;
					out<=202;
				end
				if(in == 149) begin
					state<=22;
					out<=203;
				end
				if(in == 150) begin
					state<=22;
					out<=204;
				end
				if(in == 151) begin
					state<=22;
					out<=205;
				end
				if(in == 152) begin
					state<=22;
					out<=206;
				end
				if(in == 153) begin
					state<=23;
					out<=207;
				end
				if(in == 154) begin
					state<=23;
					out<=208;
				end
				if(in == 155) begin
					state<=23;
					out<=209;
				end
				if(in == 156) begin
					state<=23;
					out<=210;
				end
				if(in == 157) begin
					state<=23;
					out<=211;
				end
				if(in == 158) begin
					state<=23;
					out<=212;
				end
				if(in == 159) begin
					state<=23;
					out<=213;
				end
				if(in == 160) begin
					state<=23;
					out<=214;
				end
				if(in == 161) begin
					state<=23;
					out<=215;
				end
				if(in == 162) begin
					state<=23;
					out<=216;
				end
				if(in == 163) begin
					state<=23;
					out<=217;
				end
				if(in == 164) begin
					state<=23;
					out<=218;
				end
				if(in == 165) begin
					state<=23;
					out<=219;
				end
				if(in == 166) begin
					state<=23;
					out<=220;
				end
				if(in == 167) begin
					state<=23;
					out<=221;
				end
				if(in == 168) begin
					state<=23;
					out<=222;
				end
				if(in == 169) begin
					state<=13;
					out<=223;
				end
				if(in == 170) begin
					state<=22;
					out<=224;
				end
				if(in == 171) begin
					state<=13;
					out<=225;
				end
				if(in == 172) begin
					state<=22;
					out<=226;
				end
				if(in == 173) begin
					state<=13;
					out<=227;
				end
				if(in == 174) begin
					state<=22;
					out<=228;
				end
				if(in == 175) begin
					state<=22;
					out<=229;
				end
				if(in == 176) begin
					state<=22;
					out<=230;
				end
				if(in == 177) begin
					state<=22;
					out<=231;
				end
				if(in == 178) begin
					state<=22;
					out<=232;
				end
				if(in == 179) begin
					state<=22;
					out<=233;
				end
				if(in == 180) begin
					state<=22;
					out<=234;
				end
				if(in == 181) begin
					state<=22;
					out<=235;
				end
				if(in == 182) begin
					state<=22;
					out<=236;
				end
				if(in == 183) begin
					state<=22;
					out<=237;
				end
				if(in == 184) begin
					state<=22;
					out<=238;
				end
				if(in == 185) begin
					state<=22;
					out<=239;
				end
				if(in == 186) begin
					state<=22;
					out<=240;
				end
				if(in == 187) begin
					state<=22;
					out<=241;
				end
				if(in == 188) begin
					state<=22;
					out<=242;
				end
				if(in == 189) begin
					state<=22;
					out<=243;
				end
				if(in == 190) begin
					state<=22;
					out<=244;
				end
				if(in == 191) begin
					state<=22;
					out<=245;
				end
				if(in == 192) begin
					state<=22;
					out<=246;
				end
				if(in == 193) begin
					state<=22;
					out<=247;
				end
				if(in == 194) begin
					state<=22;
					out<=248;
				end
				if(in == 195) begin
					state<=22;
					out<=249;
				end
				if(in == 196) begin
					state<=22;
					out<=250;
				end
				if(in == 197) begin
					state<=22;
					out<=251;
				end
				if(in == 198) begin
					state<=22;
					out<=252;
				end
				if(in == 199) begin
					state<=22;
					out<=253;
				end
				if(in == 200) begin
					state<=22;
					out<=254;
				end
				if(in == 201) begin
					state<=22;
					out<=255;
				end
				if(in == 202) begin
					state<=22;
					out<=0;
				end
				if(in == 203) begin
					state<=22;
					out<=1;
				end
				if(in == 204) begin
					state<=22;
					out<=2;
				end
				if(in == 205) begin
					state<=23;
					out<=3;
				end
				if(in == 206) begin
					state<=23;
					out<=4;
				end
				if(in == 207) begin
					state<=23;
					out<=5;
				end
				if(in == 208) begin
					state<=23;
					out<=6;
				end
				if(in == 209) begin
					state<=23;
					out<=7;
				end
				if(in == 210) begin
					state<=23;
					out<=8;
				end
				if(in == 211) begin
					state<=23;
					out<=9;
				end
				if(in == 212) begin
					state<=23;
					out<=10;
				end
				if(in == 213) begin
					state<=23;
					out<=11;
				end
				if(in == 214) begin
					state<=23;
					out<=12;
				end
				if(in == 215) begin
					state<=23;
					out<=13;
				end
				if(in == 216) begin
					state<=23;
					out<=14;
				end
				if(in == 217) begin
					state<=23;
					out<=15;
				end
				if(in == 218) begin
					state<=23;
					out<=16;
				end
				if(in == 219) begin
					state<=23;
					out<=17;
				end
				if(in == 220) begin
					state<=23;
					out<=18;
				end
				if(in == 221) begin
					state<=2;
					out<=19;
				end
				if(in == 222) begin
					state<=2;
					out<=20;
				end
				if(in == 223) begin
					state<=2;
					out<=21;
				end
				if(in == 224) begin
					state<=2;
					out<=22;
				end
				if(in == 225) begin
					state<=2;
					out<=23;
				end
				if(in == 226) begin
					state<=2;
					out<=24;
				end
				if(in == 227) begin
					state<=2;
					out<=25;
				end
				if(in == 228) begin
					state<=2;
					out<=26;
				end
				if(in == 229) begin
					state<=2;
					out<=27;
				end
				if(in == 230) begin
					state<=2;
					out<=28;
				end
				if(in == 231) begin
					state<=2;
					out<=29;
				end
				if(in == 232) begin
					state<=2;
					out<=30;
				end
				if(in == 233) begin
					state<=13;
					out<=31;
				end
				if(in == 234) begin
					state<=22;
					out<=32;
				end
				if(in == 235) begin
					state<=13;
					out<=33;
				end
				if(in == 236) begin
					state<=22;
					out<=34;
				end
				if(in == 237) begin
					state<=13;
					out<=35;
				end
				if(in == 238) begin
					state<=22;
					out<=36;
				end
				if(in == 239) begin
					state<=22;
					out<=37;
				end
				if(in == 240) begin
					state<=22;
					out<=38;
				end
				if(in == 241) begin
					state<=22;
					out<=39;
				end
				if(in == 242) begin
					state<=22;
					out<=40;
				end
				if(in == 243) begin
					state<=22;
					out<=41;
				end
				if(in == 244) begin
					state<=22;
					out<=42;
				end
				if(in == 245) begin
					state<=22;
					out<=43;
				end
				if(in == 246) begin
					state<=22;
					out<=44;
				end
				if(in == 247) begin
					state<=22;
					out<=45;
				end
				if(in == 248) begin
					state<=22;
					out<=46;
				end
				if(in == 249) begin
					state<=22;
					out<=47;
				end
				if(in == 250) begin
					state<=22;
					out<=48;
				end
				if(in == 251) begin
					state<=22;
					out<=49;
				end
				if(in == 252) begin
					state<=22;
					out<=50;
				end
				if(in == 253) begin
					state<=22;
					out<=51;
				end
				if(in == 254) begin
					state<=22;
					out<=52;
				end
				if(in == 255) begin
					state<=22;
					out<=53;
				end
				if(in == 256) begin
					state<=22;
					out<=54;
				end
				if(in == 257) begin
					state<=22;
					out<=55;
				end
				if(in == 258) begin
					state<=22;
					out<=56;
				end
				if(in == 259) begin
					state<=22;
					out<=57;
				end
				if(in == 260) begin
					state<=22;
					out<=58;
				end
				if(in == 261) begin
					state<=22;
					out<=59;
				end
				if(in == 262) begin
					state<=22;
					out<=60;
				end
				if(in == 263) begin
					state<=22;
					out<=61;
				end
				if(in == 264) begin
					state<=22;
					out<=62;
				end
				if(in == 265) begin
					state<=22;
					out<=63;
				end
				if(in == 266) begin
					state<=22;
					out<=64;
				end
				if(in == 267) begin
					state<=22;
					out<=65;
				end
				if(in == 268) begin
					state<=22;
					out<=66;
				end
				if(in == 269) begin
					state<=23;
					out<=67;
				end
				if(in == 270) begin
					state<=23;
					out<=68;
				end
				if(in == 271) begin
					state<=23;
					out<=69;
				end
				if(in == 272) begin
					state<=23;
					out<=70;
				end
				if(in == 273) begin
					state<=23;
					out<=71;
				end
				if(in == 274) begin
					state<=23;
					out<=72;
				end
				if(in == 275) begin
					state<=23;
					out<=73;
				end
				if(in == 276) begin
					state<=23;
					out<=74;
				end
				if(in == 277) begin
					state<=23;
					out<=75;
				end
				if(in == 278) begin
					state<=23;
					out<=76;
				end
				if(in == 279) begin
					state<=23;
					out<=77;
				end
				if(in == 280) begin
					state<=23;
					out<=78;
				end
				if(in == 281) begin
					state<=23;
					out<=79;
				end
				if(in == 282) begin
					state<=23;
					out<=80;
				end
				if(in == 283) begin
					state<=23;
					out<=81;
				end
				if(in == 284) begin
					state<=23;
					out<=82;
				end
				if(in == 285) begin
					state<=13;
					out<=83;
				end
				if(in == 286) begin
					state<=22;
					out<=84;
				end
				if(in == 287) begin
					state<=13;
					out<=85;
				end
				if(in == 288) begin
					state<=22;
					out<=86;
				end
				if(in == 289) begin
					state<=13;
					out<=87;
				end
				if(in == 290) begin
					state<=22;
					out<=88;
				end
				if(in == 291) begin
					state<=22;
					out<=89;
				end
				if(in == 292) begin
					state<=22;
					out<=90;
				end
				if(in == 293) begin
					state<=22;
					out<=91;
				end
				if(in == 294) begin
					state<=22;
					out<=92;
				end
				if(in == 295) begin
					state<=22;
					out<=93;
				end
				if(in == 296) begin
					state<=22;
					out<=94;
				end
				if(in == 297) begin
					state<=22;
					out<=95;
				end
				if(in == 298) begin
					state<=22;
					out<=96;
				end
				if(in == 299) begin
					state<=22;
					out<=97;
				end
				if(in == 300) begin
					state<=22;
					out<=98;
				end
				if(in == 301) begin
					state<=22;
					out<=99;
				end
				if(in == 302) begin
					state<=22;
					out<=100;
				end
				if(in == 303) begin
					state<=22;
					out<=101;
				end
				if(in == 304) begin
					state<=22;
					out<=102;
				end
				if(in == 305) begin
					state<=22;
					out<=103;
				end
				if(in == 306) begin
					state<=22;
					out<=104;
				end
				if(in == 307) begin
					state<=22;
					out<=105;
				end
				if(in == 308) begin
					state<=22;
					out<=106;
				end
				if(in == 309) begin
					state<=22;
					out<=107;
				end
				if(in == 310) begin
					state<=22;
					out<=108;
				end
				if(in == 311) begin
					state<=22;
					out<=109;
				end
				if(in == 312) begin
					state<=22;
					out<=110;
				end
				if(in == 313) begin
					state<=22;
					out<=111;
				end
				if(in == 314) begin
					state<=22;
					out<=112;
				end
				if(in == 315) begin
					state<=22;
					out<=113;
				end
				if(in == 316) begin
					state<=22;
					out<=114;
				end
				if(in == 317) begin
					state<=22;
					out<=115;
				end
				if(in == 318) begin
					state<=22;
					out<=116;
				end
				if(in == 319) begin
					state<=22;
					out<=117;
				end
				if(in == 320) begin
					state<=22;
					out<=118;
				end
				if(in == 321) begin
					state<=23;
					out<=119;
				end
				if(in == 322) begin
					state<=23;
					out<=120;
				end
				if(in == 323) begin
					state<=23;
					out<=121;
				end
				if(in == 324) begin
					state<=23;
					out<=122;
				end
				if(in == 325) begin
					state<=23;
					out<=123;
				end
				if(in == 326) begin
					state<=23;
					out<=124;
				end
				if(in == 327) begin
					state<=23;
					out<=125;
				end
				if(in == 328) begin
					state<=23;
					out<=126;
				end
				if(in == 329) begin
					state<=23;
					out<=127;
				end
				if(in == 330) begin
					state<=23;
					out<=128;
				end
				if(in == 331) begin
					state<=23;
					out<=129;
				end
				if(in == 332) begin
					state<=23;
					out<=130;
				end
				if(in == 333) begin
					state<=23;
					out<=131;
				end
				if(in == 334) begin
					state<=23;
					out<=132;
				end
				if(in == 335) begin
					state<=23;
					out<=133;
				end
				if(in == 336) begin
					state<=23;
					out<=134;
				end
				if(in == 337) begin
					state<=2;
					out<=135;
				end
				if(in == 338) begin
					state<=2;
					out<=136;
				end
				if(in == 339) begin
					state<=2;
					out<=137;
				end
				if(in == 340) begin
					state<=2;
					out<=138;
				end
				if(in == 341) begin
					state<=2;
					out<=139;
				end
				if(in == 342) begin
					state<=2;
					out<=140;
				end
				if(in == 343) begin
					state<=2;
					out<=141;
				end
				if(in == 344) begin
					state<=2;
					out<=142;
				end
				if(in == 345) begin
					state<=2;
					out<=143;
				end
				if(in == 346) begin
					state<=2;
					out<=144;
				end
				if(in == 347) begin
					state<=2;
					out<=145;
				end
				if(in == 348) begin
					state<=2;
					out<=146;
				end
				if(in == 349) begin
					state<=13;
					out<=147;
				end
				if(in == 350) begin
					state<=22;
					out<=148;
				end
				if(in == 351) begin
					state<=13;
					out<=149;
				end
				if(in == 352) begin
					state<=22;
					out<=150;
				end
				if(in == 353) begin
					state<=13;
					out<=151;
				end
				if(in == 354) begin
					state<=22;
					out<=152;
				end
				if(in == 355) begin
					state<=22;
					out<=153;
				end
				if(in == 356) begin
					state<=22;
					out<=154;
				end
				if(in == 357) begin
					state<=22;
					out<=155;
				end
				if(in == 358) begin
					state<=22;
					out<=156;
				end
				if(in == 359) begin
					state<=22;
					out<=157;
				end
				if(in == 360) begin
					state<=22;
					out<=158;
				end
				if(in == 361) begin
					state<=22;
					out<=159;
				end
				if(in == 362) begin
					state<=22;
					out<=160;
				end
				if(in == 363) begin
					state<=22;
					out<=161;
				end
				if(in == 364) begin
					state<=22;
					out<=162;
				end
				if(in == 365) begin
					state<=22;
					out<=163;
				end
				if(in == 366) begin
					state<=22;
					out<=164;
				end
				if(in == 367) begin
					state<=22;
					out<=165;
				end
				if(in == 368) begin
					state<=22;
					out<=166;
				end
				if(in == 369) begin
					state<=22;
					out<=167;
				end
				if(in == 370) begin
					state<=22;
					out<=168;
				end
				if(in == 371) begin
					state<=22;
					out<=169;
				end
				if(in == 372) begin
					state<=22;
					out<=170;
				end
				if(in == 373) begin
					state<=22;
					out<=171;
				end
				if(in == 374) begin
					state<=22;
					out<=172;
				end
				if(in == 375) begin
					state<=22;
					out<=173;
				end
				if(in == 376) begin
					state<=22;
					out<=174;
				end
				if(in == 377) begin
					state<=22;
					out<=175;
				end
				if(in == 378) begin
					state<=22;
					out<=176;
				end
				if(in == 379) begin
					state<=22;
					out<=177;
				end
				if(in == 380) begin
					state<=22;
					out<=178;
				end
				if(in == 381) begin
					state<=22;
					out<=179;
				end
				if(in == 382) begin
					state<=22;
					out<=180;
				end
				if(in == 383) begin
					state<=22;
					out<=181;
				end
				if(in == 384) begin
					state<=22;
					out<=182;
				end
				if(in == 385) begin
					state<=23;
					out<=183;
				end
				if(in == 386) begin
					state<=23;
					out<=184;
				end
				if(in == 387) begin
					state<=23;
					out<=185;
				end
				if(in == 388) begin
					state<=23;
					out<=186;
				end
				if(in == 389) begin
					state<=23;
					out<=187;
				end
				if(in == 390) begin
					state<=23;
					out<=188;
				end
				if(in == 391) begin
					state<=23;
					out<=189;
				end
				if(in == 392) begin
					state<=23;
					out<=190;
				end
				if(in == 393) begin
					state<=23;
					out<=191;
				end
				if(in == 394) begin
					state<=23;
					out<=192;
				end
				if(in == 395) begin
					state<=23;
					out<=193;
				end
				if(in == 396) begin
					state<=23;
					out<=194;
				end
				if(in == 397) begin
					state<=23;
					out<=195;
				end
				if(in == 398) begin
					state<=23;
					out<=196;
				end
				if(in == 399) begin
					state<=23;
					out<=197;
				end
				if(in == 400) begin
					state<=23;
					out<=198;
				end
				if(in == 401) begin
					state<=13;
					out<=199;
				end
				if(in == 402) begin
					state<=22;
					out<=200;
				end
				if(in == 403) begin
					state<=13;
					out<=201;
				end
				if(in == 404) begin
					state<=22;
					out<=202;
				end
				if(in == 405) begin
					state<=13;
					out<=203;
				end
				if(in == 406) begin
					state<=22;
					out<=204;
				end
				if(in == 407) begin
					state<=22;
					out<=205;
				end
				if(in == 408) begin
					state<=22;
					out<=206;
				end
				if(in == 409) begin
					state<=22;
					out<=207;
				end
				if(in == 410) begin
					state<=22;
					out<=208;
				end
				if(in == 411) begin
					state<=22;
					out<=209;
				end
				if(in == 412) begin
					state<=22;
					out<=210;
				end
				if(in == 413) begin
					state<=22;
					out<=211;
				end
				if(in == 414) begin
					state<=22;
					out<=212;
				end
				if(in == 415) begin
					state<=22;
					out<=213;
				end
				if(in == 416) begin
					state<=22;
					out<=214;
				end
				if(in == 417) begin
					state<=22;
					out<=215;
				end
				if(in == 418) begin
					state<=22;
					out<=216;
				end
				if(in == 419) begin
					state<=22;
					out<=217;
				end
				if(in == 420) begin
					state<=22;
					out<=218;
				end
				if(in == 421) begin
					state<=22;
					out<=219;
				end
				if(in == 422) begin
					state<=22;
					out<=220;
				end
				if(in == 423) begin
					state<=22;
					out<=221;
				end
				if(in == 424) begin
					state<=22;
					out<=222;
				end
				if(in == 425) begin
					state<=22;
					out<=223;
				end
				if(in == 426) begin
					state<=22;
					out<=224;
				end
				if(in == 427) begin
					state<=22;
					out<=225;
				end
				if(in == 428) begin
					state<=22;
					out<=226;
				end
				if(in == 429) begin
					state<=22;
					out<=227;
				end
				if(in == 430) begin
					state<=22;
					out<=228;
				end
				if(in == 431) begin
					state<=22;
					out<=229;
				end
				if(in == 432) begin
					state<=22;
					out<=230;
				end
				if(in == 433) begin
					state<=22;
					out<=231;
				end
				if(in == 434) begin
					state<=22;
					out<=232;
				end
				if(in == 435) begin
					state<=22;
					out<=233;
				end
				if(in == 436) begin
					state<=22;
					out<=234;
				end
				if(in == 437) begin
					state<=23;
					out<=235;
				end
				if(in == 438) begin
					state<=23;
					out<=236;
				end
				if(in == 439) begin
					state<=23;
					out<=237;
				end
				if(in == 440) begin
					state<=23;
					out<=238;
				end
				if(in == 441) begin
					state<=23;
					out<=239;
				end
				if(in == 442) begin
					state<=23;
					out<=240;
				end
				if(in == 443) begin
					state<=23;
					out<=241;
				end
				if(in == 444) begin
					state<=23;
					out<=242;
				end
				if(in == 445) begin
					state<=23;
					out<=243;
				end
				if(in == 446) begin
					state<=23;
					out<=244;
				end
				if(in == 447) begin
					state<=23;
					out<=245;
				end
				if(in == 448) begin
					state<=23;
					out<=246;
				end
				if(in == 449) begin
					state<=23;
					out<=247;
				end
				if(in == 450) begin
					state<=23;
					out<=248;
				end
				if(in == 451) begin
					state<=23;
					out<=249;
				end
				if(in == 452) begin
					state<=23;
					out<=250;
				end
				if(in == 453) begin
					state<=2;
					out<=251;
				end
				if(in == 454) begin
					state<=2;
					out<=252;
				end
				if(in == 455) begin
					state<=2;
					out<=253;
				end
				if(in == 456) begin
					state<=2;
					out<=254;
				end
				if(in == 457) begin
					state<=2;
					out<=255;
				end
				if(in == 458) begin
					state<=2;
					out<=0;
				end
				if(in == 459) begin
					state<=2;
					out<=1;
				end
				if(in == 460) begin
					state<=2;
					out<=2;
				end
				if(in == 461) begin
					state<=2;
					out<=3;
				end
				if(in == 462) begin
					state<=2;
					out<=4;
				end
				if(in == 463) begin
					state<=2;
					out<=5;
				end
				if(in == 464) begin
					state<=2;
					out<=6;
				end
				if(in == 465) begin
					state<=13;
					out<=7;
				end
				if(in == 466) begin
					state<=22;
					out<=8;
				end
				if(in == 467) begin
					state<=13;
					out<=9;
				end
				if(in == 468) begin
					state<=22;
					out<=10;
				end
				if(in == 469) begin
					state<=13;
					out<=11;
				end
				if(in == 470) begin
					state<=22;
					out<=12;
				end
				if(in == 471) begin
					state<=22;
					out<=13;
				end
				if(in == 472) begin
					state<=22;
					out<=14;
				end
				if(in == 473) begin
					state<=22;
					out<=15;
				end
				if(in == 474) begin
					state<=22;
					out<=16;
				end
				if(in == 475) begin
					state<=22;
					out<=17;
				end
				if(in == 476) begin
					state<=22;
					out<=18;
				end
				if(in == 477) begin
					state<=22;
					out<=19;
				end
				if(in == 478) begin
					state<=22;
					out<=20;
				end
				if(in == 479) begin
					state<=22;
					out<=21;
				end
				if(in == 480) begin
					state<=22;
					out<=22;
				end
				if(in == 481) begin
					state<=22;
					out<=23;
				end
				if(in == 482) begin
					state<=22;
					out<=24;
				end
				if(in == 483) begin
					state<=22;
					out<=25;
				end
				if(in == 484) begin
					state<=22;
					out<=26;
				end
				if(in == 485) begin
					state<=22;
					out<=27;
				end
				if(in == 486) begin
					state<=22;
					out<=28;
				end
				if(in == 487) begin
					state<=22;
					out<=29;
				end
				if(in == 488) begin
					state<=22;
					out<=30;
				end
				if(in == 489) begin
					state<=22;
					out<=31;
				end
				if(in == 490) begin
					state<=22;
					out<=32;
				end
				if(in == 491) begin
					state<=22;
					out<=33;
				end
				if(in == 492) begin
					state<=22;
					out<=34;
				end
				if(in == 493) begin
					state<=22;
					out<=35;
				end
				if(in == 494) begin
					state<=22;
					out<=36;
				end
				if(in == 495) begin
					state<=22;
					out<=37;
				end
				if(in == 496) begin
					state<=22;
					out<=38;
				end
				if(in == 497) begin
					state<=22;
					out<=39;
				end
				if(in == 498) begin
					state<=22;
					out<=40;
				end
				if(in == 499) begin
					state<=22;
					out<=41;
				end
				if(in == 500) begin
					state<=22;
					out<=42;
				end
				if(in == 501) begin
					state<=23;
					out<=43;
				end
				if(in == 502) begin
					state<=23;
					out<=44;
				end
				if(in == 503) begin
					state<=23;
					out<=45;
				end
				if(in == 504) begin
					state<=23;
					out<=46;
				end
				if(in == 505) begin
					state<=23;
					out<=47;
				end
				if(in == 506) begin
					state<=23;
					out<=48;
				end
				if(in == 507) begin
					state<=23;
					out<=49;
				end
				if(in == 508) begin
					state<=23;
					out<=50;
				end
				if(in == 509) begin
					state<=23;
					out<=51;
				end
				if(in == 510) begin
					state<=23;
					out<=52;
				end
				if(in == 511) begin
					state<=23;
					out<=53;
				end
				if(in == 512) begin
					state<=23;
					out<=54;
				end
				if(in == 513) begin
					state<=23;
					out<=55;
				end
				if(in == 514) begin
					state<=23;
					out<=56;
				end
				if(in == 515) begin
					state<=23;
					out<=57;
				end
				if(in == 516) begin
					state<=23;
					out<=58;
				end
				if(in == 517) begin
					state<=13;
					out<=59;
				end
				if(in == 518) begin
					state<=22;
					out<=60;
				end
				if(in == 519) begin
					state<=13;
					out<=61;
				end
				if(in == 520) begin
					state<=22;
					out<=62;
				end
				if(in == 521) begin
					state<=13;
					out<=63;
				end
				if(in == 522) begin
					state<=22;
					out<=64;
				end
				if(in == 523) begin
					state<=22;
					out<=65;
				end
				if(in == 524) begin
					state<=22;
					out<=66;
				end
				if(in == 525) begin
					state<=22;
					out<=67;
				end
				if(in == 526) begin
					state<=22;
					out<=68;
				end
				if(in == 527) begin
					state<=22;
					out<=69;
				end
				if(in == 528) begin
					state<=22;
					out<=70;
				end
				if(in == 529) begin
					state<=22;
					out<=71;
				end
				if(in == 530) begin
					state<=22;
					out<=72;
				end
				if(in == 531) begin
					state<=22;
					out<=73;
				end
				if(in == 532) begin
					state<=22;
					out<=74;
				end
				if(in == 533) begin
					state<=22;
					out<=75;
				end
				if(in == 534) begin
					state<=22;
					out<=76;
				end
				if(in == 535) begin
					state<=22;
					out<=77;
				end
				if(in == 536) begin
					state<=22;
					out<=78;
				end
				if(in == 537) begin
					state<=22;
					out<=79;
				end
				if(in == 538) begin
					state<=22;
					out<=80;
				end
				if(in == 539) begin
					state<=22;
					out<=81;
				end
				if(in == 540) begin
					state<=22;
					out<=82;
				end
				if(in == 541) begin
					state<=22;
					out<=83;
				end
				if(in == 542) begin
					state<=22;
					out<=84;
				end
				if(in == 543) begin
					state<=22;
					out<=85;
				end
				if(in == 544) begin
					state<=22;
					out<=86;
				end
				if(in == 545) begin
					state<=22;
					out<=87;
				end
				if(in == 546) begin
					state<=22;
					out<=88;
				end
				if(in == 547) begin
					state<=22;
					out<=89;
				end
				if(in == 548) begin
					state<=22;
					out<=90;
				end
				if(in == 549) begin
					state<=22;
					out<=91;
				end
				if(in == 550) begin
					state<=22;
					out<=92;
				end
				if(in == 551) begin
					state<=22;
					out<=93;
				end
				if(in == 552) begin
					state<=22;
					out<=94;
				end
				if(in == 553) begin
					state<=23;
					out<=95;
				end
				if(in == 554) begin
					state<=23;
					out<=96;
				end
				if(in == 555) begin
					state<=23;
					out<=97;
				end
				if(in == 556) begin
					state<=23;
					out<=98;
				end
				if(in == 557) begin
					state<=23;
					out<=99;
				end
				if(in == 558) begin
					state<=23;
					out<=100;
				end
				if(in == 559) begin
					state<=23;
					out<=101;
				end
				if(in == 560) begin
					state<=23;
					out<=102;
				end
				if(in == 561) begin
					state<=23;
					out<=103;
				end
				if(in == 562) begin
					state<=23;
					out<=104;
				end
				if(in == 563) begin
					state<=23;
					out<=105;
				end
				if(in == 564) begin
					state<=23;
					out<=106;
				end
				if(in == 565) begin
					state<=23;
					out<=107;
				end
				if(in == 566) begin
					state<=23;
					out<=108;
				end
				if(in == 567) begin
					state<=23;
					out<=109;
				end
				if(in == 568) begin
					state<=23;
					out<=110;
				end
				if(in == 569) begin
					state<=2;
					out<=111;
				end
				if(in == 570) begin
					state<=2;
					out<=112;
				end
				if(in == 571) begin
					state<=2;
					out<=113;
				end
				if(in == 572) begin
					state<=2;
					out<=114;
				end
				if(in == 573) begin
					state<=2;
					out<=115;
				end
				if(in == 574) begin
					state<=2;
					out<=116;
				end
				if(in == 575) begin
					state<=2;
					out<=117;
				end
				if(in == 576) begin
					state<=2;
					out<=118;
				end
				if(in == 577) begin
					state<=2;
					out<=119;
				end
				if(in == 578) begin
					state<=2;
					out<=120;
				end
				if(in == 579) begin
					state<=2;
					out<=121;
				end
				if(in == 580) begin
					state<=2;
					out<=122;
				end
				if(in == 581) begin
					state<=13;
					out<=123;
				end
				if(in == 582) begin
					state<=22;
					out<=124;
				end
				if(in == 583) begin
					state<=13;
					out<=125;
				end
				if(in == 584) begin
					state<=22;
					out<=126;
				end
				if(in == 585) begin
					state<=13;
					out<=127;
				end
				if(in == 586) begin
					state<=22;
					out<=128;
				end
				if(in == 587) begin
					state<=22;
					out<=129;
				end
				if(in == 588) begin
					state<=22;
					out<=130;
				end
				if(in == 589) begin
					state<=22;
					out<=131;
				end
				if(in == 590) begin
					state<=22;
					out<=132;
				end
				if(in == 591) begin
					state<=22;
					out<=133;
				end
				if(in == 592) begin
					state<=22;
					out<=134;
				end
				if(in == 593) begin
					state<=22;
					out<=135;
				end
				if(in == 594) begin
					state<=22;
					out<=136;
				end
				if(in == 595) begin
					state<=22;
					out<=137;
				end
				if(in == 596) begin
					state<=22;
					out<=138;
				end
				if(in == 597) begin
					state<=22;
					out<=139;
				end
				if(in == 598) begin
					state<=22;
					out<=140;
				end
				if(in == 599) begin
					state<=22;
					out<=141;
				end
				if(in == 600) begin
					state<=22;
					out<=142;
				end
				if(in == 601) begin
					state<=22;
					out<=143;
				end
				if(in == 602) begin
					state<=22;
					out<=144;
				end
				if(in == 603) begin
					state<=22;
					out<=145;
				end
				if(in == 604) begin
					state<=22;
					out<=146;
				end
				if(in == 605) begin
					state<=22;
					out<=147;
				end
				if(in == 606) begin
					state<=22;
					out<=148;
				end
				if(in == 607) begin
					state<=22;
					out<=149;
				end
				if(in == 608) begin
					state<=22;
					out<=150;
				end
				if(in == 609) begin
					state<=22;
					out<=151;
				end
				if(in == 610) begin
					state<=22;
					out<=152;
				end
				if(in == 611) begin
					state<=22;
					out<=153;
				end
				if(in == 612) begin
					state<=22;
					out<=154;
				end
				if(in == 613) begin
					state<=22;
					out<=155;
				end
				if(in == 614) begin
					state<=22;
					out<=156;
				end
				if(in == 615) begin
					state<=22;
					out<=157;
				end
				if(in == 616) begin
					state<=22;
					out<=158;
				end
				if(in == 617) begin
					state<=23;
					out<=159;
				end
				if(in == 618) begin
					state<=23;
					out<=160;
				end
				if(in == 619) begin
					state<=23;
					out<=161;
				end
				if(in == 620) begin
					state<=23;
					out<=162;
				end
				if(in == 621) begin
					state<=23;
					out<=163;
				end
				if(in == 622) begin
					state<=23;
					out<=164;
				end
				if(in == 623) begin
					state<=23;
					out<=165;
				end
				if(in == 624) begin
					state<=23;
					out<=166;
				end
				if(in == 625) begin
					state<=23;
					out<=167;
				end
				if(in == 626) begin
					state<=23;
					out<=168;
				end
				if(in == 627) begin
					state<=23;
					out<=169;
				end
				if(in == 628) begin
					state<=23;
					out<=170;
				end
				if(in == 629) begin
					state<=23;
					out<=171;
				end
				if(in == 630) begin
					state<=23;
					out<=172;
				end
				if(in == 631) begin
					state<=23;
					out<=173;
				end
				if(in == 632) begin
					state<=23;
					out<=174;
				end
				if(in == 633) begin
					state<=13;
					out<=175;
				end
				if(in == 634) begin
					state<=22;
					out<=176;
				end
				if(in == 635) begin
					state<=13;
					out<=177;
				end
				if(in == 636) begin
					state<=22;
					out<=178;
				end
				if(in == 637) begin
					state<=13;
					out<=179;
				end
				if(in == 638) begin
					state<=22;
					out<=180;
				end
				if(in == 639) begin
					state<=22;
					out<=181;
				end
				if(in == 640) begin
					state<=22;
					out<=182;
				end
				if(in == 641) begin
					state<=22;
					out<=183;
				end
				if(in == 642) begin
					state<=22;
					out<=184;
				end
				if(in == 643) begin
					state<=22;
					out<=185;
				end
				if(in == 644) begin
					state<=22;
					out<=186;
				end
				if(in == 645) begin
					state<=22;
					out<=187;
				end
				if(in == 646) begin
					state<=22;
					out<=188;
				end
				if(in == 647) begin
					state<=22;
					out<=189;
				end
				if(in == 648) begin
					state<=22;
					out<=190;
				end
				if(in == 649) begin
					state<=22;
					out<=191;
				end
				if(in == 650) begin
					state<=22;
					out<=192;
				end
				if(in == 651) begin
					state<=22;
					out<=193;
				end
				if(in == 652) begin
					state<=22;
					out<=194;
				end
				if(in == 653) begin
					state<=22;
					out<=195;
				end
				if(in == 654) begin
					state<=22;
					out<=196;
				end
				if(in == 655) begin
					state<=22;
					out<=197;
				end
				if(in == 656) begin
					state<=22;
					out<=198;
				end
				if(in == 657) begin
					state<=22;
					out<=199;
				end
				if(in == 658) begin
					state<=22;
					out<=200;
				end
				if(in == 659) begin
					state<=22;
					out<=201;
				end
				if(in == 660) begin
					state<=22;
					out<=202;
				end
				if(in == 661) begin
					state<=22;
					out<=203;
				end
				if(in == 662) begin
					state<=22;
					out<=204;
				end
				if(in == 663) begin
					state<=22;
					out<=205;
				end
				if(in == 664) begin
					state<=22;
					out<=206;
				end
				if(in == 665) begin
					state<=22;
					out<=207;
				end
				if(in == 666) begin
					state<=22;
					out<=208;
				end
				if(in == 667) begin
					state<=22;
					out<=209;
				end
				if(in == 668) begin
					state<=22;
					out<=210;
				end
				if(in == 669) begin
					state<=23;
					out<=211;
				end
				if(in == 670) begin
					state<=23;
					out<=212;
				end
				if(in == 671) begin
					state<=23;
					out<=213;
				end
				if(in == 672) begin
					state<=23;
					out<=214;
				end
				if(in == 673) begin
					state<=23;
					out<=215;
				end
				if(in == 674) begin
					state<=23;
					out<=216;
				end
				if(in == 675) begin
					state<=23;
					out<=217;
				end
				if(in == 676) begin
					state<=23;
					out<=218;
				end
				if(in == 677) begin
					state<=23;
					out<=219;
				end
				if(in == 678) begin
					state<=23;
					out<=220;
				end
				if(in == 679) begin
					state<=23;
					out<=221;
				end
				if(in == 680) begin
					state<=23;
					out<=222;
				end
				if(in == 681) begin
					state<=23;
					out<=223;
				end
				if(in == 682) begin
					state<=23;
					out<=224;
				end
				if(in == 683) begin
					state<=23;
					out<=225;
				end
				if(in == 684) begin
					state<=23;
					out<=226;
				end
				if(in == 685) begin
					state<=2;
					out<=227;
				end
				if(in == 686) begin
					state<=2;
					out<=228;
				end
				if(in == 687) begin
					state<=2;
					out<=229;
				end
				if(in == 688) begin
					state<=2;
					out<=230;
				end
				if(in == 689) begin
					state<=2;
					out<=231;
				end
				if(in == 690) begin
					state<=2;
					out<=232;
				end
				if(in == 691) begin
					state<=2;
					out<=233;
				end
				if(in == 692) begin
					state<=2;
					out<=234;
				end
				if(in == 693) begin
					state<=2;
					out<=235;
				end
				if(in == 694) begin
					state<=2;
					out<=236;
				end
				if(in == 695) begin
					state<=2;
					out<=237;
				end
				if(in == 696) begin
					state<=2;
					out<=238;
				end
				if(in == 697) begin
					state<=13;
					out<=239;
				end
				if(in == 698) begin
					state<=22;
					out<=240;
				end
				if(in == 699) begin
					state<=13;
					out<=241;
				end
				if(in == 700) begin
					state<=22;
					out<=242;
				end
				if(in == 701) begin
					state<=13;
					out<=243;
				end
				if(in == 702) begin
					state<=22;
					out<=244;
				end
				if(in == 703) begin
					state<=22;
					out<=245;
				end
				if(in == 704) begin
					state<=22;
					out<=246;
				end
				if(in == 705) begin
					state<=22;
					out<=247;
				end
				if(in == 706) begin
					state<=22;
					out<=248;
				end
				if(in == 707) begin
					state<=22;
					out<=249;
				end
				if(in == 708) begin
					state<=22;
					out<=250;
				end
				if(in == 709) begin
					state<=22;
					out<=251;
				end
				if(in == 710) begin
					state<=22;
					out<=252;
				end
				if(in == 711) begin
					state<=22;
					out<=253;
				end
				if(in == 712) begin
					state<=22;
					out<=254;
				end
				if(in == 713) begin
					state<=22;
					out<=255;
				end
				if(in == 714) begin
					state<=22;
					out<=0;
				end
				if(in == 715) begin
					state<=22;
					out<=1;
				end
				if(in == 716) begin
					state<=22;
					out<=2;
				end
				if(in == 717) begin
					state<=22;
					out<=3;
				end
				if(in == 718) begin
					state<=22;
					out<=4;
				end
				if(in == 719) begin
					state<=22;
					out<=5;
				end
				if(in == 720) begin
					state<=22;
					out<=6;
				end
				if(in == 721) begin
					state<=22;
					out<=7;
				end
				if(in == 722) begin
					state<=22;
					out<=8;
				end
				if(in == 723) begin
					state<=22;
					out<=9;
				end
				if(in == 724) begin
					state<=22;
					out<=10;
				end
				if(in == 725) begin
					state<=22;
					out<=11;
				end
				if(in == 726) begin
					state<=22;
					out<=12;
				end
				if(in == 727) begin
					state<=22;
					out<=13;
				end
				if(in == 728) begin
					state<=22;
					out<=14;
				end
				if(in == 729) begin
					state<=22;
					out<=15;
				end
				if(in == 730) begin
					state<=22;
					out<=16;
				end
				if(in == 731) begin
					state<=22;
					out<=17;
				end
				if(in == 732) begin
					state<=22;
					out<=18;
				end
				if(in == 733) begin
					state<=23;
					out<=19;
				end
				if(in == 734) begin
					state<=23;
					out<=20;
				end
				if(in == 735) begin
					state<=23;
					out<=21;
				end
				if(in == 736) begin
					state<=23;
					out<=22;
				end
				if(in == 737) begin
					state<=23;
					out<=23;
				end
				if(in == 738) begin
					state<=23;
					out<=24;
				end
				if(in == 739) begin
					state<=23;
					out<=25;
				end
				if(in == 740) begin
					state<=23;
					out<=26;
				end
				if(in == 741) begin
					state<=23;
					out<=27;
				end
				if(in == 742) begin
					state<=23;
					out<=28;
				end
				if(in == 743) begin
					state<=23;
					out<=29;
				end
				if(in == 744) begin
					state<=23;
					out<=30;
				end
				if(in == 745) begin
					state<=23;
					out<=31;
				end
				if(in == 746) begin
					state<=23;
					out<=32;
				end
				if(in == 747) begin
					state<=23;
					out<=33;
				end
				if(in == 748) begin
					state<=23;
					out<=34;
				end
				if(in == 749) begin
					state<=13;
					out<=35;
				end
				if(in == 750) begin
					state<=22;
					out<=36;
				end
				if(in == 751) begin
					state<=13;
					out<=37;
				end
				if(in == 752) begin
					state<=22;
					out<=38;
				end
				if(in == 753) begin
					state<=13;
					out<=39;
				end
				if(in == 754) begin
					state<=22;
					out<=40;
				end
				if(in == 755) begin
					state<=22;
					out<=41;
				end
				if(in == 756) begin
					state<=22;
					out<=42;
				end
				if(in == 757) begin
					state<=22;
					out<=43;
				end
				if(in == 758) begin
					state<=22;
					out<=44;
				end
				if(in == 759) begin
					state<=22;
					out<=45;
				end
				if(in == 760) begin
					state<=22;
					out<=46;
				end
				if(in == 761) begin
					state<=22;
					out<=47;
				end
				if(in == 762) begin
					state<=22;
					out<=48;
				end
				if(in == 763) begin
					state<=22;
					out<=49;
				end
				if(in == 764) begin
					state<=22;
					out<=50;
				end
				if(in == 765) begin
					state<=22;
					out<=51;
				end
				if(in == 766) begin
					state<=22;
					out<=52;
				end
				if(in == 767) begin
					state<=22;
					out<=53;
				end
				if(in == 768) begin
					state<=22;
					out<=54;
				end
				if(in == 769) begin
					state<=22;
					out<=55;
				end
				if(in == 770) begin
					state<=22;
					out<=56;
				end
				if(in == 771) begin
					state<=22;
					out<=57;
				end
				if(in == 772) begin
					state<=22;
					out<=58;
				end
				if(in == 773) begin
					state<=22;
					out<=59;
				end
				if(in == 774) begin
					state<=22;
					out<=60;
				end
				if(in == 775) begin
					state<=22;
					out<=61;
				end
				if(in == 776) begin
					state<=22;
					out<=62;
				end
				if(in == 777) begin
					state<=22;
					out<=63;
				end
				if(in == 778) begin
					state<=22;
					out<=64;
				end
				if(in == 779) begin
					state<=22;
					out<=65;
				end
				if(in == 780) begin
					state<=22;
					out<=66;
				end
				if(in == 781) begin
					state<=22;
					out<=67;
				end
				if(in == 782) begin
					state<=22;
					out<=68;
				end
				if(in == 783) begin
					state<=22;
					out<=69;
				end
				if(in == 784) begin
					state<=22;
					out<=70;
				end
				if(in == 785) begin
					state<=23;
					out<=71;
				end
				if(in == 786) begin
					state<=23;
					out<=72;
				end
				if(in == 787) begin
					state<=23;
					out<=73;
				end
				if(in == 788) begin
					state<=23;
					out<=74;
				end
				if(in == 789) begin
					state<=23;
					out<=75;
				end
				if(in == 790) begin
					state<=23;
					out<=76;
				end
				if(in == 791) begin
					state<=23;
					out<=77;
				end
				if(in == 792) begin
					state<=23;
					out<=78;
				end
				if(in == 793) begin
					state<=23;
					out<=79;
				end
				if(in == 794) begin
					state<=23;
					out<=80;
				end
				if(in == 795) begin
					state<=23;
					out<=81;
				end
				if(in == 796) begin
					state<=23;
					out<=82;
				end
				if(in == 797) begin
					state<=23;
					out<=83;
				end
				if(in == 798) begin
					state<=23;
					out<=84;
				end
				if(in == 799) begin
					state<=23;
					out<=85;
				end
				if(in == 800) begin
					state<=23;
					out<=86;
				end
				if(in == 801) begin
					state<=2;
					out<=87;
				end
				if(in == 802) begin
					state<=2;
					out<=88;
				end
				if(in == 803) begin
					state<=2;
					out<=89;
				end
				if(in == 804) begin
					state<=2;
					out<=90;
				end
				if(in == 805) begin
					state<=2;
					out<=91;
				end
				if(in == 806) begin
					state<=2;
					out<=92;
				end
				if(in == 807) begin
					state<=2;
					out<=93;
				end
				if(in == 808) begin
					state<=2;
					out<=94;
				end
				if(in == 809) begin
					state<=2;
					out<=95;
				end
				if(in == 810) begin
					state<=2;
					out<=96;
				end
				if(in == 811) begin
					state<=2;
					out<=97;
				end
				if(in == 812) begin
					state<=2;
					out<=98;
				end
				if(in == 813) begin
					state<=13;
					out<=99;
				end
				if(in == 814) begin
					state<=22;
					out<=100;
				end
				if(in == 815) begin
					state<=13;
					out<=101;
				end
				if(in == 816) begin
					state<=22;
					out<=102;
				end
				if(in == 817) begin
					state<=13;
					out<=103;
				end
				if(in == 818) begin
					state<=22;
					out<=104;
				end
				if(in == 819) begin
					state<=22;
					out<=105;
				end
				if(in == 820) begin
					state<=22;
					out<=106;
				end
				if(in == 821) begin
					state<=22;
					out<=107;
				end
				if(in == 822) begin
					state<=22;
					out<=108;
				end
				if(in == 823) begin
					state<=22;
					out<=109;
				end
				if(in == 824) begin
					state<=22;
					out<=110;
				end
				if(in == 825) begin
					state<=22;
					out<=111;
				end
				if(in == 826) begin
					state<=22;
					out<=112;
				end
				if(in == 827) begin
					state<=22;
					out<=113;
				end
				if(in == 828) begin
					state<=22;
					out<=114;
				end
				if(in == 829) begin
					state<=22;
					out<=115;
				end
				if(in == 830) begin
					state<=22;
					out<=116;
				end
				if(in == 831) begin
					state<=22;
					out<=117;
				end
				if(in == 832) begin
					state<=22;
					out<=118;
				end
				if(in == 833) begin
					state<=22;
					out<=119;
				end
				if(in == 834) begin
					state<=22;
					out<=120;
				end
				if(in == 835) begin
					state<=22;
					out<=121;
				end
				if(in == 836) begin
					state<=22;
					out<=122;
				end
				if(in == 837) begin
					state<=22;
					out<=123;
				end
				if(in == 838) begin
					state<=22;
					out<=124;
				end
				if(in == 839) begin
					state<=22;
					out<=125;
				end
				if(in == 840) begin
					state<=22;
					out<=126;
				end
				if(in == 841) begin
					state<=22;
					out<=127;
				end
				if(in == 842) begin
					state<=22;
					out<=128;
				end
				if(in == 843) begin
					state<=22;
					out<=129;
				end
				if(in == 844) begin
					state<=22;
					out<=130;
				end
				if(in == 845) begin
					state<=22;
					out<=131;
				end
				if(in == 846) begin
					state<=22;
					out<=132;
				end
				if(in == 847) begin
					state<=22;
					out<=133;
				end
				if(in == 848) begin
					state<=22;
					out<=134;
				end
				if(in == 849) begin
					state<=23;
					out<=135;
				end
				if(in == 850) begin
					state<=23;
					out<=136;
				end
				if(in == 851) begin
					state<=23;
					out<=137;
				end
				if(in == 852) begin
					state<=23;
					out<=138;
				end
				if(in == 853) begin
					state<=23;
					out<=139;
				end
				if(in == 854) begin
					state<=23;
					out<=140;
				end
				if(in == 855) begin
					state<=23;
					out<=141;
				end
				if(in == 856) begin
					state<=23;
					out<=142;
				end
				if(in == 857) begin
					state<=23;
					out<=143;
				end
				if(in == 858) begin
					state<=23;
					out<=144;
				end
				if(in == 859) begin
					state<=23;
					out<=145;
				end
				if(in == 860) begin
					state<=23;
					out<=146;
				end
				if(in == 861) begin
					state<=23;
					out<=147;
				end
				if(in == 862) begin
					state<=23;
					out<=148;
				end
				if(in == 863) begin
					state<=23;
					out<=149;
				end
				if(in == 864) begin
					state<=23;
					out<=150;
				end
				if(in == 865) begin
					state<=13;
					out<=151;
				end
				if(in == 866) begin
					state<=22;
					out<=152;
				end
				if(in == 867) begin
					state<=13;
					out<=153;
				end
				if(in == 868) begin
					state<=22;
					out<=154;
				end
				if(in == 869) begin
					state<=13;
					out<=155;
				end
				if(in == 870) begin
					state<=22;
					out<=156;
				end
				if(in == 871) begin
					state<=22;
					out<=157;
				end
				if(in == 872) begin
					state<=22;
					out<=158;
				end
				if(in == 873) begin
					state<=22;
					out<=159;
				end
				if(in == 874) begin
					state<=22;
					out<=160;
				end
				if(in == 875) begin
					state<=22;
					out<=161;
				end
				if(in == 876) begin
					state<=22;
					out<=162;
				end
				if(in == 877) begin
					state<=22;
					out<=163;
				end
				if(in == 878) begin
					state<=22;
					out<=164;
				end
				if(in == 879) begin
					state<=22;
					out<=165;
				end
				if(in == 880) begin
					state<=22;
					out<=166;
				end
				if(in == 881) begin
					state<=22;
					out<=167;
				end
				if(in == 882) begin
					state<=22;
					out<=168;
				end
				if(in == 883) begin
					state<=22;
					out<=169;
				end
				if(in == 884) begin
					state<=22;
					out<=170;
				end
				if(in == 885) begin
					state<=22;
					out<=171;
				end
				if(in == 886) begin
					state<=22;
					out<=172;
				end
				if(in == 887) begin
					state<=22;
					out<=173;
				end
				if(in == 888) begin
					state<=22;
					out<=174;
				end
				if(in == 889) begin
					state<=22;
					out<=175;
				end
				if(in == 890) begin
					state<=22;
					out<=176;
				end
				if(in == 891) begin
					state<=22;
					out<=177;
				end
				if(in == 892) begin
					state<=22;
					out<=178;
				end
				if(in == 893) begin
					state<=22;
					out<=179;
				end
				if(in == 894) begin
					state<=22;
					out<=180;
				end
				if(in == 895) begin
					state<=22;
					out<=181;
				end
				if(in == 896) begin
					state<=22;
					out<=182;
				end
				if(in == 897) begin
					state<=22;
					out<=183;
				end
				if(in == 898) begin
					state<=22;
					out<=184;
				end
				if(in == 899) begin
					state<=22;
					out<=185;
				end
				if(in == 900) begin
					state<=22;
					out<=186;
				end
				if(in == 901) begin
					state<=23;
					out<=187;
				end
				if(in == 902) begin
					state<=23;
					out<=188;
				end
				if(in == 903) begin
					state<=23;
					out<=189;
				end
				if(in == 904) begin
					state<=23;
					out<=190;
				end
				if(in == 905) begin
					state<=23;
					out<=191;
				end
				if(in == 906) begin
					state<=23;
					out<=192;
				end
				if(in == 907) begin
					state<=23;
					out<=193;
				end
				if(in == 908) begin
					state<=23;
					out<=194;
				end
				if(in == 909) begin
					state<=23;
					out<=195;
				end
				if(in == 910) begin
					state<=23;
					out<=196;
				end
				if(in == 911) begin
					state<=23;
					out<=197;
				end
				if(in == 912) begin
					state<=23;
					out<=198;
				end
				if(in == 913) begin
					state<=23;
					out<=199;
				end
				if(in == 914) begin
					state<=23;
					out<=200;
				end
				if(in == 915) begin
					state<=23;
					out<=201;
				end
				if(in == 916) begin
					state<=23;
					out<=202;
				end
				if(in == 917) begin
					state<=2;
					out<=203;
				end
				if(in == 918) begin
					state<=2;
					out<=204;
				end
				if(in == 919) begin
					state<=2;
					out<=205;
				end
				if(in == 920) begin
					state<=2;
					out<=206;
				end
				if(in == 921) begin
					state<=2;
					out<=207;
				end
				if(in == 922) begin
					state<=2;
					out<=208;
				end
				if(in == 923) begin
					state<=2;
					out<=209;
				end
				if(in == 924) begin
					state<=2;
					out<=210;
				end
				if(in == 925) begin
					state<=2;
					out<=211;
				end
				if(in == 926) begin
					state<=2;
					out<=212;
				end
				if(in == 927) begin
					state<=2;
					out<=213;
				end
				if(in == 928) begin
					state<=2;
					out<=214;
				end
			end
			23: begin
				if(in == 0) begin
					state<=13;
					out<=215;
				end
				if(in == 1) begin
					state<=1;
					out<=216;
				end
				if(in == 2) begin
					state<=23;
					out<=217;
				end
				if(in == 3) begin
					state<=13;
					out<=218;
				end
				if(in == 4) begin
					state<=23;
					out<=219;
				end
				if(in == 5) begin
					state<=13;
					out<=220;
				end
				if(in == 6) begin
					state<=23;
					out<=221;
				end
				if(in == 7) begin
					state<=23;
					out<=222;
				end
				if(in == 8) begin
					state<=23;
					out<=223;
				end
				if(in == 9) begin
					state<=23;
					out<=224;
				end
				if(in == 10) begin
					state<=23;
					out<=225;
				end
				if(in == 11) begin
					state<=23;
					out<=226;
				end
				if(in == 12) begin
					state<=23;
					out<=227;
				end
				if(in == 13) begin
					state<=23;
					out<=228;
				end
				if(in == 14) begin
					state<=23;
					out<=229;
				end
				if(in == 15) begin
					state<=23;
					out<=230;
				end
				if(in == 16) begin
					state<=23;
					out<=231;
				end
				if(in == 17) begin
					state<=23;
					out<=232;
				end
				if(in == 18) begin
					state<=23;
					out<=233;
				end
				if(in == 19) begin
					state<=23;
					out<=234;
				end
				if(in == 20) begin
					state<=23;
					out<=235;
				end
				if(in == 21) begin
					state<=23;
					out<=236;
				end
				if(in == 22) begin
					state<=23;
					out<=237;
				end
				if(in == 23) begin
					state<=23;
					out<=238;
				end
				if(in == 24) begin
					state<=23;
					out<=239;
				end
				if(in == 25) begin
					state<=23;
					out<=240;
				end
				if(in == 26) begin
					state<=23;
					out<=241;
				end
				if(in == 27) begin
					state<=23;
					out<=242;
				end
				if(in == 28) begin
					state<=23;
					out<=243;
				end
				if(in == 29) begin
					state<=23;
					out<=244;
				end
				if(in == 30) begin
					state<=23;
					out<=245;
				end
				if(in == 31) begin
					state<=23;
					out<=246;
				end
				if(in == 32) begin
					state<=23;
					out<=247;
				end
				if(in == 33) begin
					state<=23;
					out<=248;
				end
				if(in == 34) begin
					state<=23;
					out<=249;
				end
				if(in == 35) begin
					state<=23;
					out<=250;
				end
				if(in == 36) begin
					state<=23;
					out<=251;
				end
				if(in == 37) begin
					state<=23;
					out<=252;
				end
				if(in == 38) begin
					state<=23;
					out<=253;
				end
				if(in == 39) begin
					state<=23;
					out<=254;
				end
				if(in == 40) begin
					state<=23;
					out<=255;
				end
				if(in == 41) begin
					state<=23;
					out<=0;
				end
				if(in == 42) begin
					state<=23;
					out<=1;
				end
				if(in == 43) begin
					state<=23;
					out<=2;
				end
				if(in == 44) begin
					state<=23;
					out<=3;
				end
				if(in == 45) begin
					state<=23;
					out<=4;
				end
				if(in == 46) begin
					state<=23;
					out<=5;
				end
				if(in == 47) begin
					state<=23;
					out<=6;
				end
				if(in == 48) begin
					state<=23;
					out<=7;
				end
				if(in == 49) begin
					state<=23;
					out<=8;
				end
				if(in == 50) begin
					state<=23;
					out<=9;
				end
				if(in == 51) begin
					state<=23;
					out<=10;
				end
				if(in == 52) begin
					state<=23;
					out<=11;
				end
				if(in == 53) begin
					state<=13;
					out<=12;
				end
				if(in == 54) begin
					state<=23;
					out<=13;
				end
				if(in == 55) begin
					state<=13;
					out<=14;
				end
				if(in == 56) begin
					state<=23;
					out<=15;
				end
				if(in == 57) begin
					state<=13;
					out<=16;
				end
				if(in == 58) begin
					state<=23;
					out<=17;
				end
				if(in == 59) begin
					state<=23;
					out<=18;
				end
				if(in == 60) begin
					state<=23;
					out<=19;
				end
				if(in == 61) begin
					state<=23;
					out<=20;
				end
				if(in == 62) begin
					state<=23;
					out<=21;
				end
				if(in == 63) begin
					state<=23;
					out<=22;
				end
				if(in == 64) begin
					state<=23;
					out<=23;
				end
				if(in == 65) begin
					state<=23;
					out<=24;
				end
				if(in == 66) begin
					state<=23;
					out<=25;
				end
				if(in == 67) begin
					state<=23;
					out<=26;
				end
				if(in == 68) begin
					state<=23;
					out<=27;
				end
				if(in == 69) begin
					state<=23;
					out<=28;
				end
				if(in == 70) begin
					state<=23;
					out<=29;
				end
				if(in == 71) begin
					state<=23;
					out<=30;
				end
				if(in == 72) begin
					state<=23;
					out<=31;
				end
				if(in == 73) begin
					state<=23;
					out<=32;
				end
				if(in == 74) begin
					state<=23;
					out<=33;
				end
				if(in == 75) begin
					state<=23;
					out<=34;
				end
				if(in == 76) begin
					state<=23;
					out<=35;
				end
				if(in == 77) begin
					state<=23;
					out<=36;
				end
				if(in == 78) begin
					state<=23;
					out<=37;
				end
				if(in == 79) begin
					state<=23;
					out<=38;
				end
				if(in == 80) begin
					state<=23;
					out<=39;
				end
				if(in == 81) begin
					state<=23;
					out<=40;
				end
				if(in == 82) begin
					state<=23;
					out<=41;
				end
				if(in == 83) begin
					state<=23;
					out<=42;
				end
				if(in == 84) begin
					state<=23;
					out<=43;
				end
				if(in == 85) begin
					state<=23;
					out<=44;
				end
				if(in == 86) begin
					state<=23;
					out<=45;
				end
				if(in == 87) begin
					state<=23;
					out<=46;
				end
				if(in == 88) begin
					state<=23;
					out<=47;
				end
				if(in == 89) begin
					state<=23;
					out<=48;
				end
				if(in == 90) begin
					state<=23;
					out<=49;
				end
				if(in == 91) begin
					state<=23;
					out<=50;
				end
				if(in == 92) begin
					state<=23;
					out<=51;
				end
				if(in == 93) begin
					state<=23;
					out<=52;
				end
				if(in == 94) begin
					state<=23;
					out<=53;
				end
				if(in == 95) begin
					state<=23;
					out<=54;
				end
				if(in == 96) begin
					state<=23;
					out<=55;
				end
				if(in == 97) begin
					state<=23;
					out<=56;
				end
				if(in == 98) begin
					state<=23;
					out<=57;
				end
				if(in == 99) begin
					state<=23;
					out<=58;
				end
				if(in == 100) begin
					state<=23;
					out<=59;
				end
				if(in == 101) begin
					state<=23;
					out<=60;
				end
				if(in == 102) begin
					state<=23;
					out<=61;
				end
				if(in == 103) begin
					state<=23;
					out<=62;
				end
				if(in == 104) begin
					state<=23;
					out<=63;
				end
				if(in == 105) begin
					state<=2;
					out<=64;
				end
				if(in == 106) begin
					state<=2;
					out<=65;
				end
				if(in == 107) begin
					state<=2;
					out<=66;
				end
				if(in == 108) begin
					state<=2;
					out<=67;
				end
				if(in == 109) begin
					state<=2;
					out<=68;
				end
				if(in == 110) begin
					state<=2;
					out<=69;
				end
				if(in == 111) begin
					state<=2;
					out<=70;
				end
				if(in == 112) begin
					state<=2;
					out<=71;
				end
				if(in == 113) begin
					state<=2;
					out<=72;
				end
				if(in == 114) begin
					state<=2;
					out<=73;
				end
				if(in == 115) begin
					state<=2;
					out<=74;
				end
				if(in == 116) begin
					state<=2;
					out<=75;
				end
				if(in == 117) begin
					state<=13;
					out<=76;
				end
				if(in == 118) begin
					state<=23;
					out<=77;
				end
				if(in == 119) begin
					state<=13;
					out<=78;
				end
				if(in == 120) begin
					state<=23;
					out<=79;
				end
				if(in == 121) begin
					state<=13;
					out<=80;
				end
				if(in == 122) begin
					state<=23;
					out<=81;
				end
				if(in == 123) begin
					state<=23;
					out<=82;
				end
				if(in == 124) begin
					state<=23;
					out<=83;
				end
				if(in == 125) begin
					state<=23;
					out<=84;
				end
				if(in == 126) begin
					state<=23;
					out<=85;
				end
				if(in == 127) begin
					state<=23;
					out<=86;
				end
				if(in == 128) begin
					state<=23;
					out<=87;
				end
				if(in == 129) begin
					state<=23;
					out<=88;
				end
				if(in == 130) begin
					state<=23;
					out<=89;
				end
				if(in == 131) begin
					state<=23;
					out<=90;
				end
				if(in == 132) begin
					state<=23;
					out<=91;
				end
				if(in == 133) begin
					state<=23;
					out<=92;
				end
				if(in == 134) begin
					state<=23;
					out<=93;
				end
				if(in == 135) begin
					state<=23;
					out<=94;
				end
				if(in == 136) begin
					state<=23;
					out<=95;
				end
				if(in == 137) begin
					state<=23;
					out<=96;
				end
				if(in == 138) begin
					state<=23;
					out<=97;
				end
				if(in == 139) begin
					state<=23;
					out<=98;
				end
				if(in == 140) begin
					state<=23;
					out<=99;
				end
				if(in == 141) begin
					state<=23;
					out<=100;
				end
				if(in == 142) begin
					state<=23;
					out<=101;
				end
				if(in == 143) begin
					state<=23;
					out<=102;
				end
				if(in == 144) begin
					state<=23;
					out<=103;
				end
				if(in == 145) begin
					state<=23;
					out<=104;
				end
				if(in == 146) begin
					state<=23;
					out<=105;
				end
				if(in == 147) begin
					state<=23;
					out<=106;
				end
				if(in == 148) begin
					state<=23;
					out<=107;
				end
				if(in == 149) begin
					state<=23;
					out<=108;
				end
				if(in == 150) begin
					state<=23;
					out<=109;
				end
				if(in == 151) begin
					state<=23;
					out<=110;
				end
				if(in == 152) begin
					state<=23;
					out<=111;
				end
				if(in == 153) begin
					state<=23;
					out<=112;
				end
				if(in == 154) begin
					state<=23;
					out<=113;
				end
				if(in == 155) begin
					state<=23;
					out<=114;
				end
				if(in == 156) begin
					state<=23;
					out<=115;
				end
				if(in == 157) begin
					state<=23;
					out<=116;
				end
				if(in == 158) begin
					state<=23;
					out<=117;
				end
				if(in == 159) begin
					state<=23;
					out<=118;
				end
				if(in == 160) begin
					state<=23;
					out<=119;
				end
				if(in == 161) begin
					state<=23;
					out<=120;
				end
				if(in == 162) begin
					state<=23;
					out<=121;
				end
				if(in == 163) begin
					state<=23;
					out<=122;
				end
				if(in == 164) begin
					state<=23;
					out<=123;
				end
				if(in == 165) begin
					state<=23;
					out<=124;
				end
				if(in == 166) begin
					state<=23;
					out<=125;
				end
				if(in == 167) begin
					state<=23;
					out<=126;
				end
				if(in == 168) begin
					state<=23;
					out<=127;
				end
				if(in == 169) begin
					state<=13;
					out<=128;
				end
				if(in == 170) begin
					state<=23;
					out<=129;
				end
				if(in == 171) begin
					state<=13;
					out<=130;
				end
				if(in == 172) begin
					state<=23;
					out<=131;
				end
				if(in == 173) begin
					state<=13;
					out<=132;
				end
				if(in == 174) begin
					state<=23;
					out<=133;
				end
				if(in == 175) begin
					state<=23;
					out<=134;
				end
				if(in == 176) begin
					state<=23;
					out<=135;
				end
				if(in == 177) begin
					state<=23;
					out<=136;
				end
				if(in == 178) begin
					state<=23;
					out<=137;
				end
				if(in == 179) begin
					state<=23;
					out<=138;
				end
				if(in == 180) begin
					state<=23;
					out<=139;
				end
				if(in == 181) begin
					state<=23;
					out<=140;
				end
				if(in == 182) begin
					state<=23;
					out<=141;
				end
				if(in == 183) begin
					state<=23;
					out<=142;
				end
				if(in == 184) begin
					state<=23;
					out<=143;
				end
				if(in == 185) begin
					state<=23;
					out<=144;
				end
				if(in == 186) begin
					state<=23;
					out<=145;
				end
				if(in == 187) begin
					state<=23;
					out<=146;
				end
				if(in == 188) begin
					state<=23;
					out<=147;
				end
				if(in == 189) begin
					state<=23;
					out<=148;
				end
				if(in == 190) begin
					state<=23;
					out<=149;
				end
				if(in == 191) begin
					state<=23;
					out<=150;
				end
				if(in == 192) begin
					state<=23;
					out<=151;
				end
				if(in == 193) begin
					state<=23;
					out<=152;
				end
				if(in == 194) begin
					state<=23;
					out<=153;
				end
				if(in == 195) begin
					state<=23;
					out<=154;
				end
				if(in == 196) begin
					state<=23;
					out<=155;
				end
				if(in == 197) begin
					state<=23;
					out<=156;
				end
				if(in == 198) begin
					state<=23;
					out<=157;
				end
				if(in == 199) begin
					state<=23;
					out<=158;
				end
				if(in == 200) begin
					state<=23;
					out<=159;
				end
				if(in == 201) begin
					state<=23;
					out<=160;
				end
				if(in == 202) begin
					state<=23;
					out<=161;
				end
				if(in == 203) begin
					state<=23;
					out<=162;
				end
				if(in == 204) begin
					state<=23;
					out<=163;
				end
				if(in == 205) begin
					state<=23;
					out<=164;
				end
				if(in == 206) begin
					state<=23;
					out<=165;
				end
				if(in == 207) begin
					state<=23;
					out<=166;
				end
				if(in == 208) begin
					state<=23;
					out<=167;
				end
				if(in == 209) begin
					state<=23;
					out<=168;
				end
				if(in == 210) begin
					state<=23;
					out<=169;
				end
				if(in == 211) begin
					state<=23;
					out<=170;
				end
				if(in == 212) begin
					state<=23;
					out<=171;
				end
				if(in == 213) begin
					state<=23;
					out<=172;
				end
				if(in == 214) begin
					state<=23;
					out<=173;
				end
				if(in == 215) begin
					state<=23;
					out<=174;
				end
				if(in == 216) begin
					state<=23;
					out<=175;
				end
				if(in == 217) begin
					state<=23;
					out<=176;
				end
				if(in == 218) begin
					state<=23;
					out<=177;
				end
				if(in == 219) begin
					state<=23;
					out<=178;
				end
				if(in == 220) begin
					state<=23;
					out<=179;
				end
				if(in == 221) begin
					state<=2;
					out<=180;
				end
				if(in == 222) begin
					state<=2;
					out<=181;
				end
				if(in == 223) begin
					state<=2;
					out<=182;
				end
				if(in == 224) begin
					state<=2;
					out<=183;
				end
				if(in == 225) begin
					state<=2;
					out<=184;
				end
				if(in == 226) begin
					state<=2;
					out<=185;
				end
				if(in == 227) begin
					state<=2;
					out<=186;
				end
				if(in == 228) begin
					state<=2;
					out<=187;
				end
				if(in == 229) begin
					state<=2;
					out<=188;
				end
				if(in == 230) begin
					state<=2;
					out<=189;
				end
				if(in == 231) begin
					state<=2;
					out<=190;
				end
				if(in == 232) begin
					state<=2;
					out<=191;
				end
				if(in == 233) begin
					state<=13;
					out<=192;
				end
				if(in == 234) begin
					state<=23;
					out<=193;
				end
				if(in == 235) begin
					state<=13;
					out<=194;
				end
				if(in == 236) begin
					state<=23;
					out<=195;
				end
				if(in == 237) begin
					state<=13;
					out<=196;
				end
				if(in == 238) begin
					state<=23;
					out<=197;
				end
				if(in == 239) begin
					state<=23;
					out<=198;
				end
				if(in == 240) begin
					state<=23;
					out<=199;
				end
				if(in == 241) begin
					state<=23;
					out<=200;
				end
				if(in == 242) begin
					state<=23;
					out<=201;
				end
				if(in == 243) begin
					state<=23;
					out<=202;
				end
				if(in == 244) begin
					state<=23;
					out<=203;
				end
				if(in == 245) begin
					state<=23;
					out<=204;
				end
				if(in == 246) begin
					state<=23;
					out<=205;
				end
				if(in == 247) begin
					state<=23;
					out<=206;
				end
				if(in == 248) begin
					state<=23;
					out<=207;
				end
				if(in == 249) begin
					state<=23;
					out<=208;
				end
				if(in == 250) begin
					state<=23;
					out<=209;
				end
				if(in == 251) begin
					state<=23;
					out<=210;
				end
				if(in == 252) begin
					state<=23;
					out<=211;
				end
				if(in == 253) begin
					state<=23;
					out<=212;
				end
				if(in == 254) begin
					state<=23;
					out<=213;
				end
				if(in == 255) begin
					state<=23;
					out<=214;
				end
				if(in == 256) begin
					state<=23;
					out<=215;
				end
				if(in == 257) begin
					state<=23;
					out<=216;
				end
				if(in == 258) begin
					state<=23;
					out<=217;
				end
				if(in == 259) begin
					state<=23;
					out<=218;
				end
				if(in == 260) begin
					state<=23;
					out<=219;
				end
				if(in == 261) begin
					state<=23;
					out<=220;
				end
				if(in == 262) begin
					state<=23;
					out<=221;
				end
				if(in == 263) begin
					state<=23;
					out<=222;
				end
				if(in == 264) begin
					state<=23;
					out<=223;
				end
				if(in == 265) begin
					state<=23;
					out<=224;
				end
				if(in == 266) begin
					state<=23;
					out<=225;
				end
				if(in == 267) begin
					state<=23;
					out<=226;
				end
				if(in == 268) begin
					state<=23;
					out<=227;
				end
				if(in == 269) begin
					state<=23;
					out<=228;
				end
				if(in == 270) begin
					state<=23;
					out<=229;
				end
				if(in == 271) begin
					state<=23;
					out<=230;
				end
				if(in == 272) begin
					state<=23;
					out<=231;
				end
				if(in == 273) begin
					state<=23;
					out<=232;
				end
				if(in == 274) begin
					state<=23;
					out<=233;
				end
				if(in == 275) begin
					state<=23;
					out<=234;
				end
				if(in == 276) begin
					state<=23;
					out<=235;
				end
				if(in == 277) begin
					state<=23;
					out<=236;
				end
				if(in == 278) begin
					state<=23;
					out<=237;
				end
				if(in == 279) begin
					state<=23;
					out<=238;
				end
				if(in == 280) begin
					state<=23;
					out<=239;
				end
				if(in == 281) begin
					state<=23;
					out<=240;
				end
				if(in == 282) begin
					state<=23;
					out<=241;
				end
				if(in == 283) begin
					state<=23;
					out<=242;
				end
				if(in == 284) begin
					state<=23;
					out<=243;
				end
				if(in == 285) begin
					state<=13;
					out<=244;
				end
				if(in == 286) begin
					state<=23;
					out<=245;
				end
				if(in == 287) begin
					state<=13;
					out<=246;
				end
				if(in == 288) begin
					state<=23;
					out<=247;
				end
				if(in == 289) begin
					state<=13;
					out<=248;
				end
				if(in == 290) begin
					state<=23;
					out<=249;
				end
				if(in == 291) begin
					state<=23;
					out<=250;
				end
				if(in == 292) begin
					state<=23;
					out<=251;
				end
				if(in == 293) begin
					state<=23;
					out<=252;
				end
				if(in == 294) begin
					state<=23;
					out<=253;
				end
				if(in == 295) begin
					state<=23;
					out<=254;
				end
				if(in == 296) begin
					state<=23;
					out<=255;
				end
				if(in == 297) begin
					state<=23;
					out<=0;
				end
				if(in == 298) begin
					state<=23;
					out<=1;
				end
				if(in == 299) begin
					state<=23;
					out<=2;
				end
				if(in == 300) begin
					state<=23;
					out<=3;
				end
				if(in == 301) begin
					state<=23;
					out<=4;
				end
				if(in == 302) begin
					state<=23;
					out<=5;
				end
				if(in == 303) begin
					state<=23;
					out<=6;
				end
				if(in == 304) begin
					state<=23;
					out<=7;
				end
				if(in == 305) begin
					state<=23;
					out<=8;
				end
				if(in == 306) begin
					state<=23;
					out<=9;
				end
				if(in == 307) begin
					state<=23;
					out<=10;
				end
				if(in == 308) begin
					state<=23;
					out<=11;
				end
				if(in == 309) begin
					state<=23;
					out<=12;
				end
				if(in == 310) begin
					state<=23;
					out<=13;
				end
				if(in == 311) begin
					state<=23;
					out<=14;
				end
				if(in == 312) begin
					state<=23;
					out<=15;
				end
				if(in == 313) begin
					state<=23;
					out<=16;
				end
				if(in == 314) begin
					state<=23;
					out<=17;
				end
				if(in == 315) begin
					state<=23;
					out<=18;
				end
				if(in == 316) begin
					state<=23;
					out<=19;
				end
				if(in == 317) begin
					state<=23;
					out<=20;
				end
				if(in == 318) begin
					state<=23;
					out<=21;
				end
				if(in == 319) begin
					state<=23;
					out<=22;
				end
				if(in == 320) begin
					state<=23;
					out<=23;
				end
				if(in == 321) begin
					state<=23;
					out<=24;
				end
				if(in == 322) begin
					state<=23;
					out<=25;
				end
				if(in == 323) begin
					state<=23;
					out<=26;
				end
				if(in == 324) begin
					state<=23;
					out<=27;
				end
				if(in == 325) begin
					state<=23;
					out<=28;
				end
				if(in == 326) begin
					state<=23;
					out<=29;
				end
				if(in == 327) begin
					state<=23;
					out<=30;
				end
				if(in == 328) begin
					state<=23;
					out<=31;
				end
				if(in == 329) begin
					state<=23;
					out<=32;
				end
				if(in == 330) begin
					state<=23;
					out<=33;
				end
				if(in == 331) begin
					state<=23;
					out<=34;
				end
				if(in == 332) begin
					state<=23;
					out<=35;
				end
				if(in == 333) begin
					state<=23;
					out<=36;
				end
				if(in == 334) begin
					state<=23;
					out<=37;
				end
				if(in == 335) begin
					state<=23;
					out<=38;
				end
				if(in == 336) begin
					state<=23;
					out<=39;
				end
				if(in == 337) begin
					state<=2;
					out<=40;
				end
				if(in == 338) begin
					state<=2;
					out<=41;
				end
				if(in == 339) begin
					state<=2;
					out<=42;
				end
				if(in == 340) begin
					state<=2;
					out<=43;
				end
				if(in == 341) begin
					state<=2;
					out<=44;
				end
				if(in == 342) begin
					state<=2;
					out<=45;
				end
				if(in == 343) begin
					state<=2;
					out<=46;
				end
				if(in == 344) begin
					state<=2;
					out<=47;
				end
				if(in == 345) begin
					state<=2;
					out<=48;
				end
				if(in == 346) begin
					state<=2;
					out<=49;
				end
				if(in == 347) begin
					state<=2;
					out<=50;
				end
				if(in == 348) begin
					state<=2;
					out<=51;
				end
				if(in == 349) begin
					state<=13;
					out<=52;
				end
				if(in == 350) begin
					state<=23;
					out<=53;
				end
				if(in == 351) begin
					state<=13;
					out<=54;
				end
				if(in == 352) begin
					state<=23;
					out<=55;
				end
				if(in == 353) begin
					state<=13;
					out<=56;
				end
				if(in == 354) begin
					state<=23;
					out<=57;
				end
				if(in == 355) begin
					state<=23;
					out<=58;
				end
				if(in == 356) begin
					state<=23;
					out<=59;
				end
				if(in == 357) begin
					state<=23;
					out<=60;
				end
				if(in == 358) begin
					state<=23;
					out<=61;
				end
				if(in == 359) begin
					state<=23;
					out<=62;
				end
				if(in == 360) begin
					state<=23;
					out<=63;
				end
				if(in == 361) begin
					state<=23;
					out<=64;
				end
				if(in == 362) begin
					state<=23;
					out<=65;
				end
				if(in == 363) begin
					state<=23;
					out<=66;
				end
				if(in == 364) begin
					state<=23;
					out<=67;
				end
				if(in == 365) begin
					state<=23;
					out<=68;
				end
				if(in == 366) begin
					state<=23;
					out<=69;
				end
				if(in == 367) begin
					state<=23;
					out<=70;
				end
				if(in == 368) begin
					state<=23;
					out<=71;
				end
				if(in == 369) begin
					state<=23;
					out<=72;
				end
				if(in == 370) begin
					state<=23;
					out<=73;
				end
				if(in == 371) begin
					state<=23;
					out<=74;
				end
				if(in == 372) begin
					state<=23;
					out<=75;
				end
				if(in == 373) begin
					state<=23;
					out<=76;
				end
				if(in == 374) begin
					state<=23;
					out<=77;
				end
				if(in == 375) begin
					state<=23;
					out<=78;
				end
				if(in == 376) begin
					state<=23;
					out<=79;
				end
				if(in == 377) begin
					state<=23;
					out<=80;
				end
				if(in == 378) begin
					state<=23;
					out<=81;
				end
				if(in == 379) begin
					state<=23;
					out<=82;
				end
				if(in == 380) begin
					state<=23;
					out<=83;
				end
				if(in == 381) begin
					state<=23;
					out<=84;
				end
				if(in == 382) begin
					state<=23;
					out<=85;
				end
				if(in == 383) begin
					state<=23;
					out<=86;
				end
				if(in == 384) begin
					state<=23;
					out<=87;
				end
				if(in == 385) begin
					state<=23;
					out<=88;
				end
				if(in == 386) begin
					state<=23;
					out<=89;
				end
				if(in == 387) begin
					state<=23;
					out<=90;
				end
				if(in == 388) begin
					state<=23;
					out<=91;
				end
				if(in == 389) begin
					state<=23;
					out<=92;
				end
				if(in == 390) begin
					state<=23;
					out<=93;
				end
				if(in == 391) begin
					state<=23;
					out<=94;
				end
				if(in == 392) begin
					state<=23;
					out<=95;
				end
				if(in == 393) begin
					state<=23;
					out<=96;
				end
				if(in == 394) begin
					state<=23;
					out<=97;
				end
				if(in == 395) begin
					state<=23;
					out<=98;
				end
				if(in == 396) begin
					state<=23;
					out<=99;
				end
				if(in == 397) begin
					state<=23;
					out<=100;
				end
				if(in == 398) begin
					state<=23;
					out<=101;
				end
				if(in == 399) begin
					state<=23;
					out<=102;
				end
				if(in == 400) begin
					state<=23;
					out<=103;
				end
				if(in == 401) begin
					state<=13;
					out<=104;
				end
				if(in == 402) begin
					state<=23;
					out<=105;
				end
				if(in == 403) begin
					state<=13;
					out<=106;
				end
				if(in == 404) begin
					state<=23;
					out<=107;
				end
				if(in == 405) begin
					state<=13;
					out<=108;
				end
				if(in == 406) begin
					state<=23;
					out<=109;
				end
				if(in == 407) begin
					state<=23;
					out<=110;
				end
				if(in == 408) begin
					state<=23;
					out<=111;
				end
				if(in == 409) begin
					state<=23;
					out<=112;
				end
				if(in == 410) begin
					state<=23;
					out<=113;
				end
				if(in == 411) begin
					state<=23;
					out<=114;
				end
				if(in == 412) begin
					state<=23;
					out<=115;
				end
				if(in == 413) begin
					state<=23;
					out<=116;
				end
				if(in == 414) begin
					state<=23;
					out<=117;
				end
				if(in == 415) begin
					state<=23;
					out<=118;
				end
				if(in == 416) begin
					state<=23;
					out<=119;
				end
				if(in == 417) begin
					state<=23;
					out<=120;
				end
				if(in == 418) begin
					state<=23;
					out<=121;
				end
				if(in == 419) begin
					state<=23;
					out<=122;
				end
				if(in == 420) begin
					state<=23;
					out<=123;
				end
				if(in == 421) begin
					state<=23;
					out<=124;
				end
				if(in == 422) begin
					state<=23;
					out<=125;
				end
				if(in == 423) begin
					state<=23;
					out<=126;
				end
				if(in == 424) begin
					state<=23;
					out<=127;
				end
				if(in == 425) begin
					state<=23;
					out<=128;
				end
				if(in == 426) begin
					state<=23;
					out<=129;
				end
				if(in == 427) begin
					state<=23;
					out<=130;
				end
				if(in == 428) begin
					state<=23;
					out<=131;
				end
				if(in == 429) begin
					state<=23;
					out<=132;
				end
				if(in == 430) begin
					state<=23;
					out<=133;
				end
				if(in == 431) begin
					state<=23;
					out<=134;
				end
				if(in == 432) begin
					state<=23;
					out<=135;
				end
				if(in == 433) begin
					state<=23;
					out<=136;
				end
				if(in == 434) begin
					state<=23;
					out<=137;
				end
				if(in == 435) begin
					state<=23;
					out<=138;
				end
				if(in == 436) begin
					state<=23;
					out<=139;
				end
				if(in == 437) begin
					state<=23;
					out<=140;
				end
				if(in == 438) begin
					state<=23;
					out<=141;
				end
				if(in == 439) begin
					state<=23;
					out<=142;
				end
				if(in == 440) begin
					state<=23;
					out<=143;
				end
				if(in == 441) begin
					state<=23;
					out<=144;
				end
				if(in == 442) begin
					state<=23;
					out<=145;
				end
				if(in == 443) begin
					state<=23;
					out<=146;
				end
				if(in == 444) begin
					state<=23;
					out<=147;
				end
				if(in == 445) begin
					state<=23;
					out<=148;
				end
				if(in == 446) begin
					state<=23;
					out<=149;
				end
				if(in == 447) begin
					state<=23;
					out<=150;
				end
				if(in == 448) begin
					state<=23;
					out<=151;
				end
				if(in == 449) begin
					state<=23;
					out<=152;
				end
				if(in == 450) begin
					state<=23;
					out<=153;
				end
				if(in == 451) begin
					state<=23;
					out<=154;
				end
				if(in == 452) begin
					state<=23;
					out<=155;
				end
				if(in == 453) begin
					state<=2;
					out<=156;
				end
				if(in == 454) begin
					state<=2;
					out<=157;
				end
				if(in == 455) begin
					state<=2;
					out<=158;
				end
				if(in == 456) begin
					state<=2;
					out<=159;
				end
				if(in == 457) begin
					state<=2;
					out<=160;
				end
				if(in == 458) begin
					state<=2;
					out<=161;
				end
				if(in == 459) begin
					state<=2;
					out<=162;
				end
				if(in == 460) begin
					state<=2;
					out<=163;
				end
				if(in == 461) begin
					state<=2;
					out<=164;
				end
				if(in == 462) begin
					state<=2;
					out<=165;
				end
				if(in == 463) begin
					state<=2;
					out<=166;
				end
				if(in == 464) begin
					state<=2;
					out<=167;
				end
				if(in == 465) begin
					state<=13;
					out<=168;
				end
				if(in == 466) begin
					state<=23;
					out<=169;
				end
				if(in == 467) begin
					state<=13;
					out<=170;
				end
				if(in == 468) begin
					state<=23;
					out<=171;
				end
				if(in == 469) begin
					state<=13;
					out<=172;
				end
				if(in == 470) begin
					state<=23;
					out<=173;
				end
				if(in == 471) begin
					state<=23;
					out<=174;
				end
				if(in == 472) begin
					state<=23;
					out<=175;
				end
				if(in == 473) begin
					state<=23;
					out<=176;
				end
				if(in == 474) begin
					state<=23;
					out<=177;
				end
				if(in == 475) begin
					state<=23;
					out<=178;
				end
				if(in == 476) begin
					state<=23;
					out<=179;
				end
				if(in == 477) begin
					state<=23;
					out<=180;
				end
				if(in == 478) begin
					state<=23;
					out<=181;
				end
				if(in == 479) begin
					state<=23;
					out<=182;
				end
				if(in == 480) begin
					state<=23;
					out<=183;
				end
				if(in == 481) begin
					state<=23;
					out<=184;
				end
				if(in == 482) begin
					state<=23;
					out<=185;
				end
				if(in == 483) begin
					state<=23;
					out<=186;
				end
				if(in == 484) begin
					state<=23;
					out<=187;
				end
				if(in == 485) begin
					state<=23;
					out<=188;
				end
				if(in == 486) begin
					state<=23;
					out<=189;
				end
				if(in == 487) begin
					state<=23;
					out<=190;
				end
				if(in == 488) begin
					state<=23;
					out<=191;
				end
				if(in == 489) begin
					state<=23;
					out<=192;
				end
				if(in == 490) begin
					state<=23;
					out<=193;
				end
				if(in == 491) begin
					state<=23;
					out<=194;
				end
				if(in == 492) begin
					state<=23;
					out<=195;
				end
				if(in == 493) begin
					state<=23;
					out<=196;
				end
				if(in == 494) begin
					state<=23;
					out<=197;
				end
				if(in == 495) begin
					state<=23;
					out<=198;
				end
				if(in == 496) begin
					state<=23;
					out<=199;
				end
				if(in == 497) begin
					state<=23;
					out<=200;
				end
				if(in == 498) begin
					state<=23;
					out<=201;
				end
				if(in == 499) begin
					state<=23;
					out<=202;
				end
				if(in == 500) begin
					state<=23;
					out<=203;
				end
				if(in == 501) begin
					state<=23;
					out<=204;
				end
				if(in == 502) begin
					state<=23;
					out<=205;
				end
				if(in == 503) begin
					state<=23;
					out<=206;
				end
				if(in == 504) begin
					state<=23;
					out<=207;
				end
				if(in == 505) begin
					state<=23;
					out<=208;
				end
				if(in == 506) begin
					state<=23;
					out<=209;
				end
				if(in == 507) begin
					state<=23;
					out<=210;
				end
				if(in == 508) begin
					state<=23;
					out<=211;
				end
				if(in == 509) begin
					state<=23;
					out<=212;
				end
				if(in == 510) begin
					state<=23;
					out<=213;
				end
				if(in == 511) begin
					state<=23;
					out<=214;
				end
				if(in == 512) begin
					state<=23;
					out<=215;
				end
				if(in == 513) begin
					state<=23;
					out<=216;
				end
				if(in == 514) begin
					state<=23;
					out<=217;
				end
				if(in == 515) begin
					state<=23;
					out<=218;
				end
				if(in == 516) begin
					state<=23;
					out<=219;
				end
				if(in == 517) begin
					state<=13;
					out<=220;
				end
				if(in == 518) begin
					state<=23;
					out<=221;
				end
				if(in == 519) begin
					state<=13;
					out<=222;
				end
				if(in == 520) begin
					state<=23;
					out<=223;
				end
				if(in == 521) begin
					state<=13;
					out<=224;
				end
				if(in == 522) begin
					state<=23;
					out<=225;
				end
				if(in == 523) begin
					state<=23;
					out<=226;
				end
				if(in == 524) begin
					state<=23;
					out<=227;
				end
				if(in == 525) begin
					state<=23;
					out<=228;
				end
				if(in == 526) begin
					state<=23;
					out<=229;
				end
				if(in == 527) begin
					state<=23;
					out<=230;
				end
				if(in == 528) begin
					state<=23;
					out<=231;
				end
				if(in == 529) begin
					state<=23;
					out<=232;
				end
				if(in == 530) begin
					state<=23;
					out<=233;
				end
				if(in == 531) begin
					state<=23;
					out<=234;
				end
				if(in == 532) begin
					state<=23;
					out<=235;
				end
				if(in == 533) begin
					state<=23;
					out<=236;
				end
				if(in == 534) begin
					state<=23;
					out<=237;
				end
				if(in == 535) begin
					state<=23;
					out<=238;
				end
				if(in == 536) begin
					state<=23;
					out<=239;
				end
				if(in == 537) begin
					state<=23;
					out<=240;
				end
				if(in == 538) begin
					state<=23;
					out<=241;
				end
				if(in == 539) begin
					state<=23;
					out<=242;
				end
				if(in == 540) begin
					state<=23;
					out<=243;
				end
				if(in == 541) begin
					state<=23;
					out<=244;
				end
				if(in == 542) begin
					state<=23;
					out<=245;
				end
				if(in == 543) begin
					state<=23;
					out<=246;
				end
				if(in == 544) begin
					state<=23;
					out<=247;
				end
				if(in == 545) begin
					state<=23;
					out<=248;
				end
				if(in == 546) begin
					state<=23;
					out<=249;
				end
				if(in == 547) begin
					state<=23;
					out<=250;
				end
				if(in == 548) begin
					state<=23;
					out<=251;
				end
				if(in == 549) begin
					state<=23;
					out<=252;
				end
				if(in == 550) begin
					state<=23;
					out<=253;
				end
				if(in == 551) begin
					state<=23;
					out<=254;
				end
				if(in == 552) begin
					state<=23;
					out<=255;
				end
				if(in == 553) begin
					state<=23;
					out<=0;
				end
				if(in == 554) begin
					state<=23;
					out<=1;
				end
				if(in == 555) begin
					state<=23;
					out<=2;
				end
				if(in == 556) begin
					state<=23;
					out<=3;
				end
				if(in == 557) begin
					state<=23;
					out<=4;
				end
				if(in == 558) begin
					state<=23;
					out<=5;
				end
				if(in == 559) begin
					state<=23;
					out<=6;
				end
				if(in == 560) begin
					state<=23;
					out<=7;
				end
				if(in == 561) begin
					state<=23;
					out<=8;
				end
				if(in == 562) begin
					state<=23;
					out<=9;
				end
				if(in == 563) begin
					state<=23;
					out<=10;
				end
				if(in == 564) begin
					state<=23;
					out<=11;
				end
				if(in == 565) begin
					state<=23;
					out<=12;
				end
				if(in == 566) begin
					state<=23;
					out<=13;
				end
				if(in == 567) begin
					state<=23;
					out<=14;
				end
				if(in == 568) begin
					state<=23;
					out<=15;
				end
				if(in == 569) begin
					state<=2;
					out<=16;
				end
				if(in == 570) begin
					state<=2;
					out<=17;
				end
				if(in == 571) begin
					state<=2;
					out<=18;
				end
				if(in == 572) begin
					state<=2;
					out<=19;
				end
				if(in == 573) begin
					state<=2;
					out<=20;
				end
				if(in == 574) begin
					state<=2;
					out<=21;
				end
				if(in == 575) begin
					state<=2;
					out<=22;
				end
				if(in == 576) begin
					state<=2;
					out<=23;
				end
				if(in == 577) begin
					state<=2;
					out<=24;
				end
				if(in == 578) begin
					state<=2;
					out<=25;
				end
				if(in == 579) begin
					state<=2;
					out<=26;
				end
				if(in == 580) begin
					state<=2;
					out<=27;
				end
				if(in == 581) begin
					state<=13;
					out<=28;
				end
				if(in == 582) begin
					state<=23;
					out<=29;
				end
				if(in == 583) begin
					state<=13;
					out<=30;
				end
				if(in == 584) begin
					state<=23;
					out<=31;
				end
				if(in == 585) begin
					state<=13;
					out<=32;
				end
				if(in == 586) begin
					state<=23;
					out<=33;
				end
				if(in == 587) begin
					state<=23;
					out<=34;
				end
				if(in == 588) begin
					state<=23;
					out<=35;
				end
				if(in == 589) begin
					state<=23;
					out<=36;
				end
				if(in == 590) begin
					state<=23;
					out<=37;
				end
				if(in == 591) begin
					state<=23;
					out<=38;
				end
				if(in == 592) begin
					state<=23;
					out<=39;
				end
				if(in == 593) begin
					state<=23;
					out<=40;
				end
				if(in == 594) begin
					state<=23;
					out<=41;
				end
				if(in == 595) begin
					state<=23;
					out<=42;
				end
				if(in == 596) begin
					state<=23;
					out<=43;
				end
				if(in == 597) begin
					state<=23;
					out<=44;
				end
				if(in == 598) begin
					state<=23;
					out<=45;
				end
				if(in == 599) begin
					state<=23;
					out<=46;
				end
				if(in == 600) begin
					state<=23;
					out<=47;
				end
				if(in == 601) begin
					state<=23;
					out<=48;
				end
				if(in == 602) begin
					state<=23;
					out<=49;
				end
				if(in == 603) begin
					state<=23;
					out<=50;
				end
				if(in == 604) begin
					state<=23;
					out<=51;
				end
				if(in == 605) begin
					state<=23;
					out<=52;
				end
				if(in == 606) begin
					state<=23;
					out<=53;
				end
				if(in == 607) begin
					state<=23;
					out<=54;
				end
				if(in == 608) begin
					state<=23;
					out<=55;
				end
				if(in == 609) begin
					state<=23;
					out<=56;
				end
				if(in == 610) begin
					state<=23;
					out<=57;
				end
				if(in == 611) begin
					state<=23;
					out<=58;
				end
				if(in == 612) begin
					state<=23;
					out<=59;
				end
				if(in == 613) begin
					state<=23;
					out<=60;
				end
				if(in == 614) begin
					state<=23;
					out<=61;
				end
				if(in == 615) begin
					state<=23;
					out<=62;
				end
				if(in == 616) begin
					state<=23;
					out<=63;
				end
				if(in == 617) begin
					state<=23;
					out<=64;
				end
				if(in == 618) begin
					state<=23;
					out<=65;
				end
				if(in == 619) begin
					state<=23;
					out<=66;
				end
				if(in == 620) begin
					state<=23;
					out<=67;
				end
				if(in == 621) begin
					state<=23;
					out<=68;
				end
				if(in == 622) begin
					state<=23;
					out<=69;
				end
				if(in == 623) begin
					state<=23;
					out<=70;
				end
				if(in == 624) begin
					state<=23;
					out<=71;
				end
				if(in == 625) begin
					state<=23;
					out<=72;
				end
				if(in == 626) begin
					state<=23;
					out<=73;
				end
				if(in == 627) begin
					state<=23;
					out<=74;
				end
				if(in == 628) begin
					state<=23;
					out<=75;
				end
				if(in == 629) begin
					state<=23;
					out<=76;
				end
				if(in == 630) begin
					state<=23;
					out<=77;
				end
				if(in == 631) begin
					state<=23;
					out<=78;
				end
				if(in == 632) begin
					state<=23;
					out<=79;
				end
				if(in == 633) begin
					state<=13;
					out<=80;
				end
				if(in == 634) begin
					state<=23;
					out<=81;
				end
				if(in == 635) begin
					state<=13;
					out<=82;
				end
				if(in == 636) begin
					state<=23;
					out<=83;
				end
				if(in == 637) begin
					state<=13;
					out<=84;
				end
				if(in == 638) begin
					state<=23;
					out<=85;
				end
				if(in == 639) begin
					state<=23;
					out<=86;
				end
				if(in == 640) begin
					state<=23;
					out<=87;
				end
				if(in == 641) begin
					state<=23;
					out<=88;
				end
				if(in == 642) begin
					state<=23;
					out<=89;
				end
				if(in == 643) begin
					state<=23;
					out<=90;
				end
				if(in == 644) begin
					state<=23;
					out<=91;
				end
				if(in == 645) begin
					state<=23;
					out<=92;
				end
				if(in == 646) begin
					state<=23;
					out<=93;
				end
				if(in == 647) begin
					state<=23;
					out<=94;
				end
				if(in == 648) begin
					state<=23;
					out<=95;
				end
				if(in == 649) begin
					state<=23;
					out<=96;
				end
				if(in == 650) begin
					state<=23;
					out<=97;
				end
				if(in == 651) begin
					state<=23;
					out<=98;
				end
				if(in == 652) begin
					state<=23;
					out<=99;
				end
				if(in == 653) begin
					state<=23;
					out<=100;
				end
				if(in == 654) begin
					state<=23;
					out<=101;
				end
				if(in == 655) begin
					state<=23;
					out<=102;
				end
				if(in == 656) begin
					state<=23;
					out<=103;
				end
				if(in == 657) begin
					state<=23;
					out<=104;
				end
				if(in == 658) begin
					state<=23;
					out<=105;
				end
				if(in == 659) begin
					state<=23;
					out<=106;
				end
				if(in == 660) begin
					state<=23;
					out<=107;
				end
				if(in == 661) begin
					state<=23;
					out<=108;
				end
				if(in == 662) begin
					state<=23;
					out<=109;
				end
				if(in == 663) begin
					state<=23;
					out<=110;
				end
				if(in == 664) begin
					state<=23;
					out<=111;
				end
				if(in == 665) begin
					state<=23;
					out<=112;
				end
				if(in == 666) begin
					state<=23;
					out<=113;
				end
				if(in == 667) begin
					state<=23;
					out<=114;
				end
				if(in == 668) begin
					state<=23;
					out<=115;
				end
				if(in == 669) begin
					state<=23;
					out<=116;
				end
				if(in == 670) begin
					state<=23;
					out<=117;
				end
				if(in == 671) begin
					state<=23;
					out<=118;
				end
				if(in == 672) begin
					state<=23;
					out<=119;
				end
				if(in == 673) begin
					state<=23;
					out<=120;
				end
				if(in == 674) begin
					state<=23;
					out<=121;
				end
				if(in == 675) begin
					state<=23;
					out<=122;
				end
				if(in == 676) begin
					state<=23;
					out<=123;
				end
				if(in == 677) begin
					state<=23;
					out<=124;
				end
				if(in == 678) begin
					state<=23;
					out<=125;
				end
				if(in == 679) begin
					state<=23;
					out<=126;
				end
				if(in == 680) begin
					state<=23;
					out<=127;
				end
				if(in == 681) begin
					state<=23;
					out<=128;
				end
				if(in == 682) begin
					state<=23;
					out<=129;
				end
				if(in == 683) begin
					state<=23;
					out<=130;
				end
				if(in == 684) begin
					state<=23;
					out<=131;
				end
				if(in == 685) begin
					state<=2;
					out<=132;
				end
				if(in == 686) begin
					state<=2;
					out<=133;
				end
				if(in == 687) begin
					state<=2;
					out<=134;
				end
				if(in == 688) begin
					state<=2;
					out<=135;
				end
				if(in == 689) begin
					state<=2;
					out<=136;
				end
				if(in == 690) begin
					state<=2;
					out<=137;
				end
				if(in == 691) begin
					state<=2;
					out<=138;
				end
				if(in == 692) begin
					state<=2;
					out<=139;
				end
				if(in == 693) begin
					state<=2;
					out<=140;
				end
				if(in == 694) begin
					state<=2;
					out<=141;
				end
				if(in == 695) begin
					state<=2;
					out<=142;
				end
				if(in == 696) begin
					state<=2;
					out<=143;
				end
				if(in == 697) begin
					state<=13;
					out<=144;
				end
				if(in == 698) begin
					state<=23;
					out<=145;
				end
				if(in == 699) begin
					state<=13;
					out<=146;
				end
				if(in == 700) begin
					state<=23;
					out<=147;
				end
				if(in == 701) begin
					state<=13;
					out<=148;
				end
				if(in == 702) begin
					state<=23;
					out<=149;
				end
				if(in == 703) begin
					state<=23;
					out<=150;
				end
				if(in == 704) begin
					state<=23;
					out<=151;
				end
				if(in == 705) begin
					state<=23;
					out<=152;
				end
				if(in == 706) begin
					state<=23;
					out<=153;
				end
				if(in == 707) begin
					state<=23;
					out<=154;
				end
				if(in == 708) begin
					state<=23;
					out<=155;
				end
				if(in == 709) begin
					state<=23;
					out<=156;
				end
				if(in == 710) begin
					state<=23;
					out<=157;
				end
				if(in == 711) begin
					state<=23;
					out<=158;
				end
				if(in == 712) begin
					state<=23;
					out<=159;
				end
				if(in == 713) begin
					state<=23;
					out<=160;
				end
				if(in == 714) begin
					state<=23;
					out<=161;
				end
				if(in == 715) begin
					state<=23;
					out<=162;
				end
				if(in == 716) begin
					state<=23;
					out<=163;
				end
				if(in == 717) begin
					state<=23;
					out<=164;
				end
				if(in == 718) begin
					state<=23;
					out<=165;
				end
				if(in == 719) begin
					state<=23;
					out<=166;
				end
				if(in == 720) begin
					state<=23;
					out<=167;
				end
				if(in == 721) begin
					state<=23;
					out<=168;
				end
				if(in == 722) begin
					state<=23;
					out<=169;
				end
				if(in == 723) begin
					state<=23;
					out<=170;
				end
				if(in == 724) begin
					state<=23;
					out<=171;
				end
				if(in == 725) begin
					state<=23;
					out<=172;
				end
				if(in == 726) begin
					state<=23;
					out<=173;
				end
				if(in == 727) begin
					state<=23;
					out<=174;
				end
				if(in == 728) begin
					state<=23;
					out<=175;
				end
				if(in == 729) begin
					state<=23;
					out<=176;
				end
				if(in == 730) begin
					state<=23;
					out<=177;
				end
				if(in == 731) begin
					state<=23;
					out<=178;
				end
				if(in == 732) begin
					state<=23;
					out<=179;
				end
				if(in == 733) begin
					state<=23;
					out<=180;
				end
				if(in == 734) begin
					state<=23;
					out<=181;
				end
				if(in == 735) begin
					state<=23;
					out<=182;
				end
				if(in == 736) begin
					state<=23;
					out<=183;
				end
				if(in == 737) begin
					state<=23;
					out<=184;
				end
				if(in == 738) begin
					state<=23;
					out<=185;
				end
				if(in == 739) begin
					state<=23;
					out<=186;
				end
				if(in == 740) begin
					state<=23;
					out<=187;
				end
				if(in == 741) begin
					state<=23;
					out<=188;
				end
				if(in == 742) begin
					state<=23;
					out<=189;
				end
				if(in == 743) begin
					state<=23;
					out<=190;
				end
				if(in == 744) begin
					state<=23;
					out<=191;
				end
				if(in == 745) begin
					state<=23;
					out<=192;
				end
				if(in == 746) begin
					state<=23;
					out<=193;
				end
				if(in == 747) begin
					state<=23;
					out<=194;
				end
				if(in == 748) begin
					state<=23;
					out<=195;
				end
				if(in == 749) begin
					state<=13;
					out<=196;
				end
				if(in == 750) begin
					state<=23;
					out<=197;
				end
				if(in == 751) begin
					state<=13;
					out<=198;
				end
				if(in == 752) begin
					state<=23;
					out<=199;
				end
				if(in == 753) begin
					state<=13;
					out<=200;
				end
				if(in == 754) begin
					state<=23;
					out<=201;
				end
				if(in == 755) begin
					state<=23;
					out<=202;
				end
				if(in == 756) begin
					state<=23;
					out<=203;
				end
				if(in == 757) begin
					state<=23;
					out<=204;
				end
				if(in == 758) begin
					state<=23;
					out<=205;
				end
				if(in == 759) begin
					state<=23;
					out<=206;
				end
				if(in == 760) begin
					state<=23;
					out<=207;
				end
				if(in == 761) begin
					state<=23;
					out<=208;
				end
				if(in == 762) begin
					state<=23;
					out<=209;
				end
				if(in == 763) begin
					state<=23;
					out<=210;
				end
				if(in == 764) begin
					state<=23;
					out<=211;
				end
				if(in == 765) begin
					state<=23;
					out<=212;
				end
				if(in == 766) begin
					state<=23;
					out<=213;
				end
				if(in == 767) begin
					state<=23;
					out<=214;
				end
				if(in == 768) begin
					state<=23;
					out<=215;
				end
				if(in == 769) begin
					state<=23;
					out<=216;
				end
				if(in == 770) begin
					state<=23;
					out<=217;
				end
				if(in == 771) begin
					state<=23;
					out<=218;
				end
				if(in == 772) begin
					state<=23;
					out<=219;
				end
				if(in == 773) begin
					state<=23;
					out<=220;
				end
				if(in == 774) begin
					state<=23;
					out<=221;
				end
				if(in == 775) begin
					state<=23;
					out<=222;
				end
				if(in == 776) begin
					state<=23;
					out<=223;
				end
				if(in == 777) begin
					state<=23;
					out<=224;
				end
				if(in == 778) begin
					state<=23;
					out<=225;
				end
				if(in == 779) begin
					state<=23;
					out<=226;
				end
				if(in == 780) begin
					state<=23;
					out<=227;
				end
				if(in == 781) begin
					state<=23;
					out<=228;
				end
				if(in == 782) begin
					state<=23;
					out<=229;
				end
				if(in == 783) begin
					state<=23;
					out<=230;
				end
				if(in == 784) begin
					state<=23;
					out<=231;
				end
				if(in == 785) begin
					state<=23;
					out<=232;
				end
				if(in == 786) begin
					state<=23;
					out<=233;
				end
				if(in == 787) begin
					state<=23;
					out<=234;
				end
				if(in == 788) begin
					state<=23;
					out<=235;
				end
				if(in == 789) begin
					state<=23;
					out<=236;
				end
				if(in == 790) begin
					state<=23;
					out<=237;
				end
				if(in == 791) begin
					state<=23;
					out<=238;
				end
				if(in == 792) begin
					state<=23;
					out<=239;
				end
				if(in == 793) begin
					state<=23;
					out<=240;
				end
				if(in == 794) begin
					state<=23;
					out<=241;
				end
				if(in == 795) begin
					state<=23;
					out<=242;
				end
				if(in == 796) begin
					state<=23;
					out<=243;
				end
				if(in == 797) begin
					state<=23;
					out<=244;
				end
				if(in == 798) begin
					state<=23;
					out<=245;
				end
				if(in == 799) begin
					state<=23;
					out<=246;
				end
				if(in == 800) begin
					state<=23;
					out<=247;
				end
				if(in == 801) begin
					state<=2;
					out<=248;
				end
				if(in == 802) begin
					state<=2;
					out<=249;
				end
				if(in == 803) begin
					state<=2;
					out<=250;
				end
				if(in == 804) begin
					state<=2;
					out<=251;
				end
				if(in == 805) begin
					state<=2;
					out<=252;
				end
				if(in == 806) begin
					state<=2;
					out<=253;
				end
				if(in == 807) begin
					state<=2;
					out<=254;
				end
				if(in == 808) begin
					state<=2;
					out<=255;
				end
				if(in == 809) begin
					state<=2;
					out<=0;
				end
				if(in == 810) begin
					state<=2;
					out<=1;
				end
				if(in == 811) begin
					state<=2;
					out<=2;
				end
				if(in == 812) begin
					state<=2;
					out<=3;
				end
				if(in == 813) begin
					state<=13;
					out<=4;
				end
				if(in == 814) begin
					state<=23;
					out<=5;
				end
				if(in == 815) begin
					state<=13;
					out<=6;
				end
				if(in == 816) begin
					state<=23;
					out<=7;
				end
				if(in == 817) begin
					state<=13;
					out<=8;
				end
				if(in == 818) begin
					state<=23;
					out<=9;
				end
				if(in == 819) begin
					state<=23;
					out<=10;
				end
				if(in == 820) begin
					state<=23;
					out<=11;
				end
				if(in == 821) begin
					state<=23;
					out<=12;
				end
				if(in == 822) begin
					state<=23;
					out<=13;
				end
				if(in == 823) begin
					state<=23;
					out<=14;
				end
				if(in == 824) begin
					state<=23;
					out<=15;
				end
				if(in == 825) begin
					state<=23;
					out<=16;
				end
				if(in == 826) begin
					state<=23;
					out<=17;
				end
				if(in == 827) begin
					state<=23;
					out<=18;
				end
				if(in == 828) begin
					state<=23;
					out<=19;
				end
				if(in == 829) begin
					state<=23;
					out<=20;
				end
				if(in == 830) begin
					state<=23;
					out<=21;
				end
				if(in == 831) begin
					state<=23;
					out<=22;
				end
				if(in == 832) begin
					state<=23;
					out<=23;
				end
				if(in == 833) begin
					state<=23;
					out<=24;
				end
				if(in == 834) begin
					state<=23;
					out<=25;
				end
				if(in == 835) begin
					state<=23;
					out<=26;
				end
				if(in == 836) begin
					state<=23;
					out<=27;
				end
				if(in == 837) begin
					state<=23;
					out<=28;
				end
				if(in == 838) begin
					state<=23;
					out<=29;
				end
				if(in == 839) begin
					state<=23;
					out<=30;
				end
				if(in == 840) begin
					state<=23;
					out<=31;
				end
				if(in == 841) begin
					state<=23;
					out<=32;
				end
				if(in == 842) begin
					state<=23;
					out<=33;
				end
				if(in == 843) begin
					state<=23;
					out<=34;
				end
				if(in == 844) begin
					state<=23;
					out<=35;
				end
				if(in == 845) begin
					state<=23;
					out<=36;
				end
				if(in == 846) begin
					state<=23;
					out<=37;
				end
				if(in == 847) begin
					state<=23;
					out<=38;
				end
				if(in == 848) begin
					state<=23;
					out<=39;
				end
				if(in == 849) begin
					state<=23;
					out<=40;
				end
				if(in == 850) begin
					state<=23;
					out<=41;
				end
				if(in == 851) begin
					state<=23;
					out<=42;
				end
				if(in == 852) begin
					state<=23;
					out<=43;
				end
				if(in == 853) begin
					state<=23;
					out<=44;
				end
				if(in == 854) begin
					state<=23;
					out<=45;
				end
				if(in == 855) begin
					state<=23;
					out<=46;
				end
				if(in == 856) begin
					state<=23;
					out<=47;
				end
				if(in == 857) begin
					state<=23;
					out<=48;
				end
				if(in == 858) begin
					state<=23;
					out<=49;
				end
				if(in == 859) begin
					state<=23;
					out<=50;
				end
				if(in == 860) begin
					state<=23;
					out<=51;
				end
				if(in == 861) begin
					state<=23;
					out<=52;
				end
				if(in == 862) begin
					state<=23;
					out<=53;
				end
				if(in == 863) begin
					state<=23;
					out<=54;
				end
				if(in == 864) begin
					state<=23;
					out<=55;
				end
				if(in == 865) begin
					state<=13;
					out<=56;
				end
				if(in == 866) begin
					state<=23;
					out<=57;
				end
				if(in == 867) begin
					state<=13;
					out<=58;
				end
				if(in == 868) begin
					state<=23;
					out<=59;
				end
				if(in == 869) begin
					state<=13;
					out<=60;
				end
				if(in == 870) begin
					state<=23;
					out<=61;
				end
				if(in == 871) begin
					state<=23;
					out<=62;
				end
				if(in == 872) begin
					state<=23;
					out<=63;
				end
				if(in == 873) begin
					state<=23;
					out<=64;
				end
				if(in == 874) begin
					state<=23;
					out<=65;
				end
				if(in == 875) begin
					state<=23;
					out<=66;
				end
				if(in == 876) begin
					state<=23;
					out<=67;
				end
				if(in == 877) begin
					state<=23;
					out<=68;
				end
				if(in == 878) begin
					state<=23;
					out<=69;
				end
				if(in == 879) begin
					state<=23;
					out<=70;
				end
				if(in == 880) begin
					state<=23;
					out<=71;
				end
				if(in == 881) begin
					state<=23;
					out<=72;
				end
				if(in == 882) begin
					state<=23;
					out<=73;
				end
				if(in == 883) begin
					state<=23;
					out<=74;
				end
				if(in == 884) begin
					state<=23;
					out<=75;
				end
				if(in == 885) begin
					state<=23;
					out<=76;
				end
				if(in == 886) begin
					state<=23;
					out<=77;
				end
				if(in == 887) begin
					state<=23;
					out<=78;
				end
				if(in == 888) begin
					state<=23;
					out<=79;
				end
				if(in == 889) begin
					state<=23;
					out<=80;
				end
				if(in == 890) begin
					state<=23;
					out<=81;
				end
				if(in == 891) begin
					state<=23;
					out<=82;
				end
				if(in == 892) begin
					state<=23;
					out<=83;
				end
				if(in == 893) begin
					state<=23;
					out<=84;
				end
				if(in == 894) begin
					state<=23;
					out<=85;
				end
				if(in == 895) begin
					state<=23;
					out<=86;
				end
				if(in == 896) begin
					state<=23;
					out<=87;
				end
				if(in == 897) begin
					state<=23;
					out<=88;
				end
				if(in == 898) begin
					state<=23;
					out<=89;
				end
				if(in == 899) begin
					state<=23;
					out<=90;
				end
				if(in == 900) begin
					state<=23;
					out<=91;
				end
				if(in == 901) begin
					state<=23;
					out<=92;
				end
				if(in == 902) begin
					state<=23;
					out<=93;
				end
				if(in == 903) begin
					state<=23;
					out<=94;
				end
				if(in == 904) begin
					state<=23;
					out<=95;
				end
				if(in == 905) begin
					state<=23;
					out<=96;
				end
				if(in == 906) begin
					state<=23;
					out<=97;
				end
				if(in == 907) begin
					state<=23;
					out<=98;
				end
				if(in == 908) begin
					state<=23;
					out<=99;
				end
				if(in == 909) begin
					state<=23;
					out<=100;
				end
				if(in == 910) begin
					state<=23;
					out<=101;
				end
				if(in == 911) begin
					state<=23;
					out<=102;
				end
				if(in == 912) begin
					state<=23;
					out<=103;
				end
				if(in == 913) begin
					state<=23;
					out<=104;
				end
				if(in == 914) begin
					state<=23;
					out<=105;
				end
				if(in == 915) begin
					state<=23;
					out<=106;
				end
				if(in == 916) begin
					state<=23;
					out<=107;
				end
				if(in == 917) begin
					state<=2;
					out<=108;
				end
				if(in == 918) begin
					state<=2;
					out<=109;
				end
				if(in == 919) begin
					state<=2;
					out<=110;
				end
				if(in == 920) begin
					state<=2;
					out<=111;
				end
				if(in == 921) begin
					state<=2;
					out<=112;
				end
				if(in == 922) begin
					state<=2;
					out<=113;
				end
				if(in == 923) begin
					state<=2;
					out<=114;
				end
				if(in == 924) begin
					state<=2;
					out<=115;
				end
				if(in == 925) begin
					state<=2;
					out<=116;
				end
				if(in == 926) begin
					state<=2;
					out<=117;
				end
				if(in == 927) begin
					state<=2;
					out<=118;
				end
				if(in == 928) begin
					state<=2;
					out<=119;
				end
			end
			24: begin
				if(in == 0) begin
					state<=24;
					out<=120;
				end
				if(in == 1) begin
					state<=1;
					out<=121;
				end
				if(in == 2) begin
					state<=24;
					out<=122;
				end
				if(in == 3) begin
					state<=24;
					out<=123;
				end
				if(in == 4) begin
					state<=24;
					out<=124;
				end
				if(in == 5) begin
					state<=24;
					out<=125;
				end
				if(in == 6) begin
					state<=24;
					out<=126;
				end
				if(in == 7) begin
					state<=24;
					out<=127;
				end
				if(in == 8) begin
					state<=24;
					out<=128;
				end
				if(in == 9) begin
					state<=24;
					out<=129;
				end
				if(in == 10) begin
					state<=24;
					out<=130;
				end
				if(in == 11) begin
					state<=24;
					out<=131;
				end
				if(in == 12) begin
					state<=24;
					out<=132;
				end
				if(in == 13) begin
					state<=24;
					out<=133;
				end
				if(in == 14) begin
					state<=24;
					out<=134;
				end
				if(in == 15) begin
					state<=24;
					out<=135;
				end
				if(in == 16) begin
					state<=24;
					out<=136;
				end
				if(in == 17) begin
					state<=24;
					out<=137;
				end
				if(in == 18) begin
					state<=24;
					out<=138;
				end
				if(in == 19) begin
					state<=24;
					out<=139;
				end
				if(in == 20) begin
					state<=24;
					out<=140;
				end
				if(in == 21) begin
					state<=24;
					out<=141;
				end
				if(in == 22) begin
					state<=24;
					out<=142;
				end
				if(in == 23) begin
					state<=24;
					out<=143;
				end
				if(in == 24) begin
					state<=24;
					out<=144;
				end
				if(in == 25) begin
					state<=24;
					out<=145;
				end
				if(in == 26) begin
					state<=24;
					out<=146;
				end
				if(in == 27) begin
					state<=24;
					out<=147;
				end
				if(in == 28) begin
					state<=24;
					out<=148;
				end
				if(in == 29) begin
					state<=24;
					out<=149;
				end
				if(in == 30) begin
					state<=24;
					out<=150;
				end
				if(in == 31) begin
					state<=24;
					out<=151;
				end
				if(in == 32) begin
					state<=24;
					out<=152;
				end
				if(in == 33) begin
					state<=24;
					out<=153;
				end
				if(in == 34) begin
					state<=24;
					out<=154;
				end
				if(in == 35) begin
					state<=24;
					out<=155;
				end
				if(in == 36) begin
					state<=24;
					out<=156;
				end
				if(in == 37) begin
					state<=24;
					out<=157;
				end
				if(in == 38) begin
					state<=24;
					out<=158;
				end
				if(in == 39) begin
					state<=24;
					out<=159;
				end
				if(in == 40) begin
					state<=24;
					out<=160;
				end
				if(in == 41) begin
					state<=24;
					out<=161;
				end
				if(in == 42) begin
					state<=24;
					out<=162;
				end
				if(in == 43) begin
					state<=24;
					out<=163;
				end
				if(in == 44) begin
					state<=24;
					out<=164;
				end
				if(in == 45) begin
					state<=24;
					out<=165;
				end
				if(in == 46) begin
					state<=24;
					out<=166;
				end
				if(in == 47) begin
					state<=24;
					out<=167;
				end
				if(in == 48) begin
					state<=24;
					out<=168;
				end
				if(in == 49) begin
					state<=24;
					out<=169;
				end
				if(in == 50) begin
					state<=24;
					out<=170;
				end
				if(in == 51) begin
					state<=24;
					out<=171;
				end
				if(in == 52) begin
					state<=24;
					out<=172;
				end
				if(in == 53) begin
					state<=24;
					out<=173;
				end
				if(in == 54) begin
					state<=24;
					out<=174;
				end
				if(in == 55) begin
					state<=24;
					out<=175;
				end
				if(in == 56) begin
					state<=24;
					out<=176;
				end
				if(in == 57) begin
					state<=24;
					out<=177;
				end
				if(in == 58) begin
					state<=24;
					out<=178;
				end
				if(in == 59) begin
					state<=24;
					out<=179;
				end
				if(in == 60) begin
					state<=24;
					out<=180;
				end
				if(in == 61) begin
					state<=24;
					out<=181;
				end
				if(in == 62) begin
					state<=24;
					out<=182;
				end
				if(in == 63) begin
					state<=24;
					out<=183;
				end
				if(in == 64) begin
					state<=24;
					out<=184;
				end
				if(in == 65) begin
					state<=24;
					out<=185;
				end
				if(in == 66) begin
					state<=24;
					out<=186;
				end
				if(in == 67) begin
					state<=24;
					out<=187;
				end
				if(in == 68) begin
					state<=24;
					out<=188;
				end
				if(in == 69) begin
					state<=24;
					out<=189;
				end
				if(in == 70) begin
					state<=24;
					out<=190;
				end
				if(in == 71) begin
					state<=24;
					out<=191;
				end
				if(in == 72) begin
					state<=24;
					out<=192;
				end
				if(in == 73) begin
					state<=24;
					out<=193;
				end
				if(in == 74) begin
					state<=24;
					out<=194;
				end
				if(in == 75) begin
					state<=24;
					out<=195;
				end
				if(in == 76) begin
					state<=24;
					out<=196;
				end
				if(in == 77) begin
					state<=24;
					out<=197;
				end
				if(in == 78) begin
					state<=24;
					out<=198;
				end
				if(in == 79) begin
					state<=24;
					out<=199;
				end
				if(in == 80) begin
					state<=24;
					out<=200;
				end
				if(in == 81) begin
					state<=24;
					out<=201;
				end
				if(in == 82) begin
					state<=24;
					out<=202;
				end
				if(in == 83) begin
					state<=24;
					out<=203;
				end
				if(in == 84) begin
					state<=24;
					out<=204;
				end
				if(in == 85) begin
					state<=24;
					out<=205;
				end
				if(in == 86) begin
					state<=24;
					out<=206;
				end
				if(in == 87) begin
					state<=24;
					out<=207;
				end
				if(in == 88) begin
					state<=24;
					out<=208;
				end
				if(in == 89) begin
					state<=24;
					out<=209;
				end
				if(in == 90) begin
					state<=24;
					out<=210;
				end
				if(in == 91) begin
					state<=24;
					out<=211;
				end
				if(in == 92) begin
					state<=24;
					out<=212;
				end
				if(in == 93) begin
					state<=24;
					out<=213;
				end
				if(in == 94) begin
					state<=24;
					out<=214;
				end
				if(in == 95) begin
					state<=24;
					out<=215;
				end
				if(in == 96) begin
					state<=24;
					out<=216;
				end
				if(in == 97) begin
					state<=24;
					out<=217;
				end
				if(in == 98) begin
					state<=24;
					out<=218;
				end
				if(in == 99) begin
					state<=24;
					out<=219;
				end
				if(in == 100) begin
					state<=24;
					out<=220;
				end
				if(in == 101) begin
					state<=24;
					out<=221;
				end
				if(in == 102) begin
					state<=24;
					out<=222;
				end
				if(in == 103) begin
					state<=24;
					out<=223;
				end
				if(in == 104) begin
					state<=24;
					out<=224;
				end
				if(in == 105) begin
					state<=24;
					out<=225;
				end
				if(in == 106) begin
					state<=24;
					out<=226;
				end
				if(in == 107) begin
					state<=24;
					out<=227;
				end
				if(in == 108) begin
					state<=24;
					out<=228;
				end
				if(in == 109) begin
					state<=24;
					out<=229;
				end
				if(in == 110) begin
					state<=24;
					out<=230;
				end
				if(in == 111) begin
					state<=24;
					out<=231;
				end
				if(in == 112) begin
					state<=24;
					out<=232;
				end
				if(in == 113) begin
					state<=24;
					out<=233;
				end
				if(in == 114) begin
					state<=24;
					out<=234;
				end
				if(in == 115) begin
					state<=24;
					out<=235;
				end
				if(in == 116) begin
					state<=24;
					out<=236;
				end
				if(in == 117) begin
					state<=24;
					out<=237;
				end
				if(in == 118) begin
					state<=24;
					out<=238;
				end
				if(in == 119) begin
					state<=24;
					out<=239;
				end
				if(in == 120) begin
					state<=24;
					out<=240;
				end
				if(in == 121) begin
					state<=24;
					out<=241;
				end
				if(in == 122) begin
					state<=24;
					out<=242;
				end
				if(in == 123) begin
					state<=24;
					out<=243;
				end
				if(in == 124) begin
					state<=24;
					out<=244;
				end
				if(in == 125) begin
					state<=24;
					out<=245;
				end
				if(in == 126) begin
					state<=24;
					out<=246;
				end
				if(in == 127) begin
					state<=24;
					out<=247;
				end
				if(in == 128) begin
					state<=24;
					out<=248;
				end
				if(in == 129) begin
					state<=24;
					out<=249;
				end
				if(in == 130) begin
					state<=24;
					out<=250;
				end
				if(in == 131) begin
					state<=24;
					out<=251;
				end
				if(in == 132) begin
					state<=24;
					out<=252;
				end
				if(in == 133) begin
					state<=24;
					out<=253;
				end
				if(in == 134) begin
					state<=24;
					out<=254;
				end
				if(in == 135) begin
					state<=24;
					out<=255;
				end
				if(in == 136) begin
					state<=24;
					out<=0;
				end
				if(in == 137) begin
					state<=24;
					out<=1;
				end
				if(in == 138) begin
					state<=24;
					out<=2;
				end
				if(in == 139) begin
					state<=24;
					out<=3;
				end
				if(in == 140) begin
					state<=24;
					out<=4;
				end
				if(in == 141) begin
					state<=24;
					out<=5;
				end
				if(in == 142) begin
					state<=24;
					out<=6;
				end
				if(in == 143) begin
					state<=24;
					out<=7;
				end
				if(in == 144) begin
					state<=24;
					out<=8;
				end
				if(in == 145) begin
					state<=24;
					out<=9;
				end
				if(in == 146) begin
					state<=24;
					out<=10;
				end
				if(in == 147) begin
					state<=24;
					out<=11;
				end
				if(in == 148) begin
					state<=24;
					out<=12;
				end
				if(in == 149) begin
					state<=24;
					out<=13;
				end
				if(in == 150) begin
					state<=24;
					out<=14;
				end
				if(in == 151) begin
					state<=24;
					out<=15;
				end
				if(in == 152) begin
					state<=24;
					out<=16;
				end
				if(in == 153) begin
					state<=24;
					out<=17;
				end
				if(in == 154) begin
					state<=24;
					out<=18;
				end
				if(in == 155) begin
					state<=24;
					out<=19;
				end
				if(in == 156) begin
					state<=24;
					out<=20;
				end
				if(in == 157) begin
					state<=24;
					out<=21;
				end
				if(in == 158) begin
					state<=24;
					out<=22;
				end
				if(in == 159) begin
					state<=24;
					out<=23;
				end
				if(in == 160) begin
					state<=24;
					out<=24;
				end
				if(in == 161) begin
					state<=24;
					out<=25;
				end
				if(in == 162) begin
					state<=24;
					out<=26;
				end
				if(in == 163) begin
					state<=24;
					out<=27;
				end
				if(in == 164) begin
					state<=24;
					out<=28;
				end
				if(in == 165) begin
					state<=24;
					out<=29;
				end
				if(in == 166) begin
					state<=24;
					out<=30;
				end
				if(in == 167) begin
					state<=24;
					out<=31;
				end
				if(in == 168) begin
					state<=24;
					out<=32;
				end
				if(in == 169) begin
					state<=24;
					out<=33;
				end
				if(in == 170) begin
					state<=24;
					out<=34;
				end
				if(in == 171) begin
					state<=24;
					out<=35;
				end
				if(in == 172) begin
					state<=24;
					out<=36;
				end
				if(in == 173) begin
					state<=24;
					out<=37;
				end
				if(in == 174) begin
					state<=24;
					out<=38;
				end
				if(in == 175) begin
					state<=24;
					out<=39;
				end
				if(in == 176) begin
					state<=24;
					out<=40;
				end
				if(in == 177) begin
					state<=24;
					out<=41;
				end
				if(in == 178) begin
					state<=24;
					out<=42;
				end
				if(in == 179) begin
					state<=24;
					out<=43;
				end
				if(in == 180) begin
					state<=24;
					out<=44;
				end
				if(in == 181) begin
					state<=24;
					out<=45;
				end
				if(in == 182) begin
					state<=24;
					out<=46;
				end
				if(in == 183) begin
					state<=24;
					out<=47;
				end
				if(in == 184) begin
					state<=24;
					out<=48;
				end
				if(in == 185) begin
					state<=24;
					out<=49;
				end
				if(in == 186) begin
					state<=24;
					out<=50;
				end
				if(in == 187) begin
					state<=24;
					out<=51;
				end
				if(in == 188) begin
					state<=24;
					out<=52;
				end
				if(in == 189) begin
					state<=24;
					out<=53;
				end
				if(in == 190) begin
					state<=24;
					out<=54;
				end
				if(in == 191) begin
					state<=24;
					out<=55;
				end
				if(in == 192) begin
					state<=24;
					out<=56;
				end
				if(in == 193) begin
					state<=24;
					out<=57;
				end
				if(in == 194) begin
					state<=24;
					out<=58;
				end
				if(in == 195) begin
					state<=24;
					out<=59;
				end
				if(in == 196) begin
					state<=24;
					out<=60;
				end
				if(in == 197) begin
					state<=24;
					out<=61;
				end
				if(in == 198) begin
					state<=24;
					out<=62;
				end
				if(in == 199) begin
					state<=24;
					out<=63;
				end
				if(in == 200) begin
					state<=24;
					out<=64;
				end
				if(in == 201) begin
					state<=24;
					out<=65;
				end
				if(in == 202) begin
					state<=24;
					out<=66;
				end
				if(in == 203) begin
					state<=24;
					out<=67;
				end
				if(in == 204) begin
					state<=24;
					out<=68;
				end
				if(in == 205) begin
					state<=24;
					out<=69;
				end
				if(in == 206) begin
					state<=24;
					out<=70;
				end
				if(in == 207) begin
					state<=24;
					out<=71;
				end
				if(in == 208) begin
					state<=24;
					out<=72;
				end
				if(in == 209) begin
					state<=24;
					out<=73;
				end
				if(in == 210) begin
					state<=24;
					out<=74;
				end
				if(in == 211) begin
					state<=24;
					out<=75;
				end
				if(in == 212) begin
					state<=24;
					out<=76;
				end
				if(in == 213) begin
					state<=24;
					out<=77;
				end
				if(in == 214) begin
					state<=24;
					out<=78;
				end
				if(in == 215) begin
					state<=24;
					out<=79;
				end
				if(in == 216) begin
					state<=24;
					out<=80;
				end
				if(in == 217) begin
					state<=24;
					out<=81;
				end
				if(in == 218) begin
					state<=24;
					out<=82;
				end
				if(in == 219) begin
					state<=24;
					out<=83;
				end
				if(in == 220) begin
					state<=24;
					out<=84;
				end
				if(in == 221) begin
					state<=24;
					out<=85;
				end
				if(in == 222) begin
					state<=24;
					out<=86;
				end
				if(in == 223) begin
					state<=24;
					out<=87;
				end
				if(in == 224) begin
					state<=24;
					out<=88;
				end
				if(in == 225) begin
					state<=24;
					out<=89;
				end
				if(in == 226) begin
					state<=24;
					out<=90;
				end
				if(in == 227) begin
					state<=24;
					out<=91;
				end
				if(in == 228) begin
					state<=24;
					out<=92;
				end
				if(in == 229) begin
					state<=24;
					out<=93;
				end
				if(in == 230) begin
					state<=24;
					out<=94;
				end
				if(in == 231) begin
					state<=24;
					out<=95;
				end
				if(in == 232) begin
					state<=24;
					out<=96;
				end
				if(in == 233) begin
					state<=24;
					out<=97;
				end
				if(in == 234) begin
					state<=24;
					out<=98;
				end
				if(in == 235) begin
					state<=24;
					out<=99;
				end
				if(in == 236) begin
					state<=24;
					out<=100;
				end
				if(in == 237) begin
					state<=24;
					out<=101;
				end
				if(in == 238) begin
					state<=24;
					out<=102;
				end
				if(in == 239) begin
					state<=24;
					out<=103;
				end
				if(in == 240) begin
					state<=24;
					out<=104;
				end
				if(in == 241) begin
					state<=24;
					out<=105;
				end
				if(in == 242) begin
					state<=24;
					out<=106;
				end
				if(in == 243) begin
					state<=24;
					out<=107;
				end
				if(in == 244) begin
					state<=24;
					out<=108;
				end
				if(in == 245) begin
					state<=24;
					out<=109;
				end
				if(in == 246) begin
					state<=24;
					out<=110;
				end
				if(in == 247) begin
					state<=24;
					out<=111;
				end
				if(in == 248) begin
					state<=24;
					out<=112;
				end
				if(in == 249) begin
					state<=24;
					out<=113;
				end
				if(in == 250) begin
					state<=24;
					out<=114;
				end
				if(in == 251) begin
					state<=24;
					out<=115;
				end
				if(in == 252) begin
					state<=24;
					out<=116;
				end
				if(in == 253) begin
					state<=24;
					out<=117;
				end
				if(in == 254) begin
					state<=24;
					out<=118;
				end
				if(in == 255) begin
					state<=24;
					out<=119;
				end
				if(in == 256) begin
					state<=24;
					out<=120;
				end
				if(in == 257) begin
					state<=24;
					out<=121;
				end
				if(in == 258) begin
					state<=24;
					out<=122;
				end
				if(in == 259) begin
					state<=24;
					out<=123;
				end
				if(in == 260) begin
					state<=24;
					out<=124;
				end
				if(in == 261) begin
					state<=24;
					out<=125;
				end
				if(in == 262) begin
					state<=24;
					out<=126;
				end
				if(in == 263) begin
					state<=24;
					out<=127;
				end
				if(in == 264) begin
					state<=24;
					out<=128;
				end
				if(in == 265) begin
					state<=24;
					out<=129;
				end
				if(in == 266) begin
					state<=24;
					out<=130;
				end
				if(in == 267) begin
					state<=24;
					out<=131;
				end
				if(in == 268) begin
					state<=24;
					out<=132;
				end
				if(in == 269) begin
					state<=24;
					out<=133;
				end
				if(in == 270) begin
					state<=24;
					out<=134;
				end
				if(in == 271) begin
					state<=24;
					out<=135;
				end
				if(in == 272) begin
					state<=24;
					out<=136;
				end
				if(in == 273) begin
					state<=24;
					out<=137;
				end
				if(in == 274) begin
					state<=24;
					out<=138;
				end
				if(in == 275) begin
					state<=24;
					out<=139;
				end
				if(in == 276) begin
					state<=24;
					out<=140;
				end
				if(in == 277) begin
					state<=24;
					out<=141;
				end
				if(in == 278) begin
					state<=24;
					out<=142;
				end
				if(in == 279) begin
					state<=24;
					out<=143;
				end
				if(in == 280) begin
					state<=24;
					out<=144;
				end
				if(in == 281) begin
					state<=24;
					out<=145;
				end
				if(in == 282) begin
					state<=24;
					out<=146;
				end
				if(in == 283) begin
					state<=24;
					out<=147;
				end
				if(in == 284) begin
					state<=24;
					out<=148;
				end
				if(in == 285) begin
					state<=24;
					out<=149;
				end
				if(in == 286) begin
					state<=24;
					out<=150;
				end
				if(in == 287) begin
					state<=24;
					out<=151;
				end
				if(in == 288) begin
					state<=24;
					out<=152;
				end
				if(in == 289) begin
					state<=24;
					out<=153;
				end
				if(in == 290) begin
					state<=24;
					out<=154;
				end
				if(in == 291) begin
					state<=24;
					out<=155;
				end
				if(in == 292) begin
					state<=24;
					out<=156;
				end
				if(in == 293) begin
					state<=24;
					out<=157;
				end
				if(in == 294) begin
					state<=24;
					out<=158;
				end
				if(in == 295) begin
					state<=24;
					out<=159;
				end
				if(in == 296) begin
					state<=24;
					out<=160;
				end
				if(in == 297) begin
					state<=24;
					out<=161;
				end
				if(in == 298) begin
					state<=24;
					out<=162;
				end
				if(in == 299) begin
					state<=24;
					out<=163;
				end
				if(in == 300) begin
					state<=24;
					out<=164;
				end
				if(in == 301) begin
					state<=24;
					out<=165;
				end
				if(in == 302) begin
					state<=24;
					out<=166;
				end
				if(in == 303) begin
					state<=24;
					out<=167;
				end
				if(in == 304) begin
					state<=24;
					out<=168;
				end
				if(in == 305) begin
					state<=24;
					out<=169;
				end
				if(in == 306) begin
					state<=24;
					out<=170;
				end
				if(in == 307) begin
					state<=24;
					out<=171;
				end
				if(in == 308) begin
					state<=24;
					out<=172;
				end
				if(in == 309) begin
					state<=24;
					out<=173;
				end
				if(in == 310) begin
					state<=24;
					out<=174;
				end
				if(in == 311) begin
					state<=24;
					out<=175;
				end
				if(in == 312) begin
					state<=24;
					out<=176;
				end
				if(in == 313) begin
					state<=24;
					out<=177;
				end
				if(in == 314) begin
					state<=24;
					out<=178;
				end
				if(in == 315) begin
					state<=24;
					out<=179;
				end
				if(in == 316) begin
					state<=24;
					out<=180;
				end
				if(in == 317) begin
					state<=24;
					out<=181;
				end
				if(in == 318) begin
					state<=24;
					out<=182;
				end
				if(in == 319) begin
					state<=24;
					out<=183;
				end
				if(in == 320) begin
					state<=24;
					out<=184;
				end
				if(in == 321) begin
					state<=24;
					out<=185;
				end
				if(in == 322) begin
					state<=24;
					out<=186;
				end
				if(in == 323) begin
					state<=24;
					out<=187;
				end
				if(in == 324) begin
					state<=24;
					out<=188;
				end
				if(in == 325) begin
					state<=24;
					out<=189;
				end
				if(in == 326) begin
					state<=24;
					out<=190;
				end
				if(in == 327) begin
					state<=24;
					out<=191;
				end
				if(in == 328) begin
					state<=24;
					out<=192;
				end
				if(in == 329) begin
					state<=24;
					out<=193;
				end
				if(in == 330) begin
					state<=24;
					out<=194;
				end
				if(in == 331) begin
					state<=24;
					out<=195;
				end
				if(in == 332) begin
					state<=24;
					out<=196;
				end
				if(in == 333) begin
					state<=24;
					out<=197;
				end
				if(in == 334) begin
					state<=24;
					out<=198;
				end
				if(in == 335) begin
					state<=24;
					out<=199;
				end
				if(in == 336) begin
					state<=24;
					out<=200;
				end
				if(in == 337) begin
					state<=24;
					out<=201;
				end
				if(in == 338) begin
					state<=24;
					out<=202;
				end
				if(in == 339) begin
					state<=24;
					out<=203;
				end
				if(in == 340) begin
					state<=24;
					out<=204;
				end
				if(in == 341) begin
					state<=24;
					out<=205;
				end
				if(in == 342) begin
					state<=24;
					out<=206;
				end
				if(in == 343) begin
					state<=24;
					out<=207;
				end
				if(in == 344) begin
					state<=24;
					out<=208;
				end
				if(in == 345) begin
					state<=24;
					out<=209;
				end
				if(in == 346) begin
					state<=24;
					out<=210;
				end
				if(in == 347) begin
					state<=24;
					out<=211;
				end
				if(in == 348) begin
					state<=24;
					out<=212;
				end
				if(in == 349) begin
					state<=24;
					out<=213;
				end
				if(in == 350) begin
					state<=24;
					out<=214;
				end
				if(in == 351) begin
					state<=24;
					out<=215;
				end
				if(in == 352) begin
					state<=24;
					out<=216;
				end
				if(in == 353) begin
					state<=24;
					out<=217;
				end
				if(in == 354) begin
					state<=24;
					out<=218;
				end
				if(in == 355) begin
					state<=24;
					out<=219;
				end
				if(in == 356) begin
					state<=24;
					out<=220;
				end
				if(in == 357) begin
					state<=24;
					out<=221;
				end
				if(in == 358) begin
					state<=24;
					out<=222;
				end
				if(in == 359) begin
					state<=24;
					out<=223;
				end
				if(in == 360) begin
					state<=24;
					out<=224;
				end
				if(in == 361) begin
					state<=24;
					out<=225;
				end
				if(in == 362) begin
					state<=24;
					out<=226;
				end
				if(in == 363) begin
					state<=24;
					out<=227;
				end
				if(in == 364) begin
					state<=24;
					out<=228;
				end
				if(in == 365) begin
					state<=24;
					out<=229;
				end
				if(in == 366) begin
					state<=24;
					out<=230;
				end
				if(in == 367) begin
					state<=24;
					out<=231;
				end
				if(in == 368) begin
					state<=24;
					out<=232;
				end
				if(in == 369) begin
					state<=24;
					out<=233;
				end
				if(in == 370) begin
					state<=24;
					out<=234;
				end
				if(in == 371) begin
					state<=24;
					out<=235;
				end
				if(in == 372) begin
					state<=24;
					out<=236;
				end
				if(in == 373) begin
					state<=24;
					out<=237;
				end
				if(in == 374) begin
					state<=24;
					out<=238;
				end
				if(in == 375) begin
					state<=24;
					out<=239;
				end
				if(in == 376) begin
					state<=24;
					out<=240;
				end
				if(in == 377) begin
					state<=24;
					out<=241;
				end
				if(in == 378) begin
					state<=24;
					out<=242;
				end
				if(in == 379) begin
					state<=24;
					out<=243;
				end
				if(in == 380) begin
					state<=24;
					out<=244;
				end
				if(in == 381) begin
					state<=24;
					out<=245;
				end
				if(in == 382) begin
					state<=24;
					out<=246;
				end
				if(in == 383) begin
					state<=24;
					out<=247;
				end
				if(in == 384) begin
					state<=24;
					out<=248;
				end
				if(in == 385) begin
					state<=24;
					out<=249;
				end
				if(in == 386) begin
					state<=24;
					out<=250;
				end
				if(in == 387) begin
					state<=24;
					out<=251;
				end
				if(in == 388) begin
					state<=24;
					out<=252;
				end
				if(in == 389) begin
					state<=24;
					out<=253;
				end
				if(in == 390) begin
					state<=24;
					out<=254;
				end
				if(in == 391) begin
					state<=24;
					out<=255;
				end
				if(in == 392) begin
					state<=24;
					out<=0;
				end
				if(in == 393) begin
					state<=24;
					out<=1;
				end
				if(in == 394) begin
					state<=24;
					out<=2;
				end
				if(in == 395) begin
					state<=24;
					out<=3;
				end
				if(in == 396) begin
					state<=24;
					out<=4;
				end
				if(in == 397) begin
					state<=24;
					out<=5;
				end
				if(in == 398) begin
					state<=24;
					out<=6;
				end
				if(in == 399) begin
					state<=24;
					out<=7;
				end
				if(in == 400) begin
					state<=24;
					out<=8;
				end
				if(in == 401) begin
					state<=24;
					out<=9;
				end
				if(in == 402) begin
					state<=24;
					out<=10;
				end
				if(in == 403) begin
					state<=24;
					out<=11;
				end
				if(in == 404) begin
					state<=24;
					out<=12;
				end
				if(in == 405) begin
					state<=24;
					out<=13;
				end
				if(in == 406) begin
					state<=24;
					out<=14;
				end
				if(in == 407) begin
					state<=24;
					out<=15;
				end
				if(in == 408) begin
					state<=24;
					out<=16;
				end
				if(in == 409) begin
					state<=24;
					out<=17;
				end
				if(in == 410) begin
					state<=24;
					out<=18;
				end
				if(in == 411) begin
					state<=24;
					out<=19;
				end
				if(in == 412) begin
					state<=24;
					out<=20;
				end
				if(in == 413) begin
					state<=24;
					out<=21;
				end
				if(in == 414) begin
					state<=24;
					out<=22;
				end
				if(in == 415) begin
					state<=24;
					out<=23;
				end
				if(in == 416) begin
					state<=24;
					out<=24;
				end
				if(in == 417) begin
					state<=24;
					out<=25;
				end
				if(in == 418) begin
					state<=24;
					out<=26;
				end
				if(in == 419) begin
					state<=24;
					out<=27;
				end
				if(in == 420) begin
					state<=24;
					out<=28;
				end
				if(in == 421) begin
					state<=24;
					out<=29;
				end
				if(in == 422) begin
					state<=24;
					out<=30;
				end
				if(in == 423) begin
					state<=24;
					out<=31;
				end
				if(in == 424) begin
					state<=24;
					out<=32;
				end
				if(in == 425) begin
					state<=24;
					out<=33;
				end
				if(in == 426) begin
					state<=24;
					out<=34;
				end
				if(in == 427) begin
					state<=24;
					out<=35;
				end
				if(in == 428) begin
					state<=24;
					out<=36;
				end
				if(in == 429) begin
					state<=24;
					out<=37;
				end
				if(in == 430) begin
					state<=24;
					out<=38;
				end
				if(in == 431) begin
					state<=24;
					out<=39;
				end
				if(in == 432) begin
					state<=24;
					out<=40;
				end
				if(in == 433) begin
					state<=24;
					out<=41;
				end
				if(in == 434) begin
					state<=24;
					out<=42;
				end
				if(in == 435) begin
					state<=24;
					out<=43;
				end
				if(in == 436) begin
					state<=24;
					out<=44;
				end
				if(in == 437) begin
					state<=24;
					out<=45;
				end
				if(in == 438) begin
					state<=24;
					out<=46;
				end
				if(in == 439) begin
					state<=24;
					out<=47;
				end
				if(in == 440) begin
					state<=24;
					out<=48;
				end
				if(in == 441) begin
					state<=24;
					out<=49;
				end
				if(in == 442) begin
					state<=24;
					out<=50;
				end
				if(in == 443) begin
					state<=24;
					out<=51;
				end
				if(in == 444) begin
					state<=24;
					out<=52;
				end
				if(in == 445) begin
					state<=24;
					out<=53;
				end
				if(in == 446) begin
					state<=24;
					out<=54;
				end
				if(in == 447) begin
					state<=24;
					out<=55;
				end
				if(in == 448) begin
					state<=24;
					out<=56;
				end
				if(in == 449) begin
					state<=24;
					out<=57;
				end
				if(in == 450) begin
					state<=24;
					out<=58;
				end
				if(in == 451) begin
					state<=24;
					out<=59;
				end
				if(in == 452) begin
					state<=24;
					out<=60;
				end
				if(in == 453) begin
					state<=24;
					out<=61;
				end
				if(in == 454) begin
					state<=24;
					out<=62;
				end
				if(in == 455) begin
					state<=24;
					out<=63;
				end
				if(in == 456) begin
					state<=24;
					out<=64;
				end
				if(in == 457) begin
					state<=24;
					out<=65;
				end
				if(in == 458) begin
					state<=24;
					out<=66;
				end
				if(in == 459) begin
					state<=24;
					out<=67;
				end
				if(in == 460) begin
					state<=24;
					out<=68;
				end
				if(in == 461) begin
					state<=24;
					out<=69;
				end
				if(in == 462) begin
					state<=24;
					out<=70;
				end
				if(in == 463) begin
					state<=24;
					out<=71;
				end
				if(in == 464) begin
					state<=24;
					out<=72;
				end
				if(in == 465) begin
					state<=1;
					out<=73;
				end
				if(in == 466) begin
					state<=1;
					out<=74;
				end
				if(in == 467) begin
					state<=1;
					out<=75;
				end
				if(in == 468) begin
					state<=1;
					out<=76;
				end
				if(in == 469) begin
					state<=1;
					out<=77;
				end
				if(in == 470) begin
					state<=1;
					out<=78;
				end
				if(in == 471) begin
					state<=1;
					out<=79;
				end
				if(in == 472) begin
					state<=1;
					out<=80;
				end
				if(in == 473) begin
					state<=1;
					out<=81;
				end
				if(in == 474) begin
					state<=1;
					out<=82;
				end
				if(in == 475) begin
					state<=1;
					out<=83;
				end
				if(in == 476) begin
					state<=1;
					out<=84;
				end
				if(in == 477) begin
					state<=1;
					out<=85;
				end
				if(in == 478) begin
					state<=1;
					out<=86;
				end
				if(in == 479) begin
					state<=1;
					out<=87;
				end
				if(in == 480) begin
					state<=1;
					out<=88;
				end
				if(in == 481) begin
					state<=1;
					out<=89;
				end
				if(in == 482) begin
					state<=1;
					out<=90;
				end
				if(in == 483) begin
					state<=1;
					out<=91;
				end
				if(in == 484) begin
					state<=1;
					out<=92;
				end
				if(in == 485) begin
					state<=1;
					out<=93;
				end
				if(in == 486) begin
					state<=1;
					out<=94;
				end
				if(in == 487) begin
					state<=1;
					out<=95;
				end
				if(in == 488) begin
					state<=1;
					out<=96;
				end
				if(in == 489) begin
					state<=1;
					out<=97;
				end
				if(in == 490) begin
					state<=1;
					out<=98;
				end
				if(in == 491) begin
					state<=1;
					out<=99;
				end
				if(in == 492) begin
					state<=1;
					out<=100;
				end
				if(in == 493) begin
					state<=1;
					out<=101;
				end
				if(in == 494) begin
					state<=1;
					out<=102;
				end
				if(in == 495) begin
					state<=1;
					out<=103;
				end
				if(in == 496) begin
					state<=1;
					out<=104;
				end
				if(in == 497) begin
					state<=1;
					out<=105;
				end
				if(in == 498) begin
					state<=1;
					out<=106;
				end
				if(in == 499) begin
					state<=1;
					out<=107;
				end
				if(in == 500) begin
					state<=1;
					out<=108;
				end
				if(in == 501) begin
					state<=1;
					out<=109;
				end
				if(in == 502) begin
					state<=1;
					out<=110;
				end
				if(in == 503) begin
					state<=1;
					out<=111;
				end
				if(in == 504) begin
					state<=1;
					out<=112;
				end
				if(in == 505) begin
					state<=1;
					out<=113;
				end
				if(in == 506) begin
					state<=1;
					out<=114;
				end
				if(in == 507) begin
					state<=1;
					out<=115;
				end
				if(in == 508) begin
					state<=1;
					out<=116;
				end
				if(in == 509) begin
					state<=1;
					out<=117;
				end
				if(in == 510) begin
					state<=1;
					out<=118;
				end
				if(in == 511) begin
					state<=1;
					out<=119;
				end
				if(in == 512) begin
					state<=1;
					out<=120;
				end
				if(in == 513) begin
					state<=1;
					out<=121;
				end
				if(in == 514) begin
					state<=1;
					out<=122;
				end
				if(in == 515) begin
					state<=1;
					out<=123;
				end
				if(in == 516) begin
					state<=1;
					out<=124;
				end
				if(in == 517) begin
					state<=1;
					out<=125;
				end
				if(in == 518) begin
					state<=1;
					out<=126;
				end
				if(in == 519) begin
					state<=1;
					out<=127;
				end
				if(in == 520) begin
					state<=1;
					out<=128;
				end
				if(in == 521) begin
					state<=1;
					out<=129;
				end
				if(in == 522) begin
					state<=1;
					out<=130;
				end
				if(in == 523) begin
					state<=1;
					out<=131;
				end
				if(in == 524) begin
					state<=1;
					out<=132;
				end
				if(in == 525) begin
					state<=1;
					out<=133;
				end
				if(in == 526) begin
					state<=1;
					out<=134;
				end
				if(in == 527) begin
					state<=1;
					out<=135;
				end
				if(in == 528) begin
					state<=1;
					out<=136;
				end
				if(in == 529) begin
					state<=1;
					out<=137;
				end
				if(in == 530) begin
					state<=1;
					out<=138;
				end
				if(in == 531) begin
					state<=1;
					out<=139;
				end
				if(in == 532) begin
					state<=1;
					out<=140;
				end
				if(in == 533) begin
					state<=1;
					out<=141;
				end
				if(in == 534) begin
					state<=1;
					out<=142;
				end
				if(in == 535) begin
					state<=1;
					out<=143;
				end
				if(in == 536) begin
					state<=1;
					out<=144;
				end
				if(in == 537) begin
					state<=1;
					out<=145;
				end
				if(in == 538) begin
					state<=1;
					out<=146;
				end
				if(in == 539) begin
					state<=1;
					out<=147;
				end
				if(in == 540) begin
					state<=1;
					out<=148;
				end
				if(in == 541) begin
					state<=1;
					out<=149;
				end
				if(in == 542) begin
					state<=1;
					out<=150;
				end
				if(in == 543) begin
					state<=1;
					out<=151;
				end
				if(in == 544) begin
					state<=1;
					out<=152;
				end
				if(in == 545) begin
					state<=1;
					out<=153;
				end
				if(in == 546) begin
					state<=1;
					out<=154;
				end
				if(in == 547) begin
					state<=1;
					out<=155;
				end
				if(in == 548) begin
					state<=1;
					out<=156;
				end
				if(in == 549) begin
					state<=1;
					out<=157;
				end
				if(in == 550) begin
					state<=1;
					out<=158;
				end
				if(in == 551) begin
					state<=1;
					out<=159;
				end
				if(in == 552) begin
					state<=1;
					out<=160;
				end
				if(in == 553) begin
					state<=1;
					out<=161;
				end
				if(in == 554) begin
					state<=1;
					out<=162;
				end
				if(in == 555) begin
					state<=1;
					out<=163;
				end
				if(in == 556) begin
					state<=1;
					out<=164;
				end
				if(in == 557) begin
					state<=1;
					out<=165;
				end
				if(in == 558) begin
					state<=1;
					out<=166;
				end
				if(in == 559) begin
					state<=1;
					out<=167;
				end
				if(in == 560) begin
					state<=1;
					out<=168;
				end
				if(in == 561) begin
					state<=1;
					out<=169;
				end
				if(in == 562) begin
					state<=1;
					out<=170;
				end
				if(in == 563) begin
					state<=1;
					out<=171;
				end
				if(in == 564) begin
					state<=1;
					out<=172;
				end
				if(in == 565) begin
					state<=1;
					out<=173;
				end
				if(in == 566) begin
					state<=1;
					out<=174;
				end
				if(in == 567) begin
					state<=1;
					out<=175;
				end
				if(in == 568) begin
					state<=1;
					out<=176;
				end
				if(in == 569) begin
					state<=1;
					out<=177;
				end
				if(in == 570) begin
					state<=1;
					out<=178;
				end
				if(in == 571) begin
					state<=1;
					out<=179;
				end
				if(in == 572) begin
					state<=1;
					out<=180;
				end
				if(in == 573) begin
					state<=1;
					out<=181;
				end
				if(in == 574) begin
					state<=1;
					out<=182;
				end
				if(in == 575) begin
					state<=1;
					out<=183;
				end
				if(in == 576) begin
					state<=1;
					out<=184;
				end
				if(in == 577) begin
					state<=1;
					out<=185;
				end
				if(in == 578) begin
					state<=1;
					out<=186;
				end
				if(in == 579) begin
					state<=1;
					out<=187;
				end
				if(in == 580) begin
					state<=1;
					out<=188;
				end
				if(in == 581) begin
					state<=1;
					out<=189;
				end
				if(in == 582) begin
					state<=1;
					out<=190;
				end
				if(in == 583) begin
					state<=1;
					out<=191;
				end
				if(in == 584) begin
					state<=1;
					out<=192;
				end
				if(in == 585) begin
					state<=1;
					out<=193;
				end
				if(in == 586) begin
					state<=1;
					out<=194;
				end
				if(in == 587) begin
					state<=1;
					out<=195;
				end
				if(in == 588) begin
					state<=1;
					out<=196;
				end
				if(in == 589) begin
					state<=1;
					out<=197;
				end
				if(in == 590) begin
					state<=1;
					out<=198;
				end
				if(in == 591) begin
					state<=1;
					out<=199;
				end
				if(in == 592) begin
					state<=1;
					out<=200;
				end
				if(in == 593) begin
					state<=1;
					out<=201;
				end
				if(in == 594) begin
					state<=1;
					out<=202;
				end
				if(in == 595) begin
					state<=1;
					out<=203;
				end
				if(in == 596) begin
					state<=1;
					out<=204;
				end
				if(in == 597) begin
					state<=1;
					out<=205;
				end
				if(in == 598) begin
					state<=1;
					out<=206;
				end
				if(in == 599) begin
					state<=1;
					out<=207;
				end
				if(in == 600) begin
					state<=1;
					out<=208;
				end
				if(in == 601) begin
					state<=1;
					out<=209;
				end
				if(in == 602) begin
					state<=1;
					out<=210;
				end
				if(in == 603) begin
					state<=1;
					out<=211;
				end
				if(in == 604) begin
					state<=1;
					out<=212;
				end
				if(in == 605) begin
					state<=1;
					out<=213;
				end
				if(in == 606) begin
					state<=1;
					out<=214;
				end
				if(in == 607) begin
					state<=1;
					out<=215;
				end
				if(in == 608) begin
					state<=1;
					out<=216;
				end
				if(in == 609) begin
					state<=1;
					out<=217;
				end
				if(in == 610) begin
					state<=1;
					out<=218;
				end
				if(in == 611) begin
					state<=1;
					out<=219;
				end
				if(in == 612) begin
					state<=1;
					out<=220;
				end
				if(in == 613) begin
					state<=1;
					out<=221;
				end
				if(in == 614) begin
					state<=1;
					out<=222;
				end
				if(in == 615) begin
					state<=1;
					out<=223;
				end
				if(in == 616) begin
					state<=1;
					out<=224;
				end
				if(in == 617) begin
					state<=1;
					out<=225;
				end
				if(in == 618) begin
					state<=1;
					out<=226;
				end
				if(in == 619) begin
					state<=1;
					out<=227;
				end
				if(in == 620) begin
					state<=1;
					out<=228;
				end
				if(in == 621) begin
					state<=1;
					out<=229;
				end
				if(in == 622) begin
					state<=1;
					out<=230;
				end
				if(in == 623) begin
					state<=1;
					out<=231;
				end
				if(in == 624) begin
					state<=1;
					out<=232;
				end
				if(in == 625) begin
					state<=1;
					out<=233;
				end
				if(in == 626) begin
					state<=1;
					out<=234;
				end
				if(in == 627) begin
					state<=1;
					out<=235;
				end
				if(in == 628) begin
					state<=1;
					out<=236;
				end
				if(in == 629) begin
					state<=1;
					out<=237;
				end
				if(in == 630) begin
					state<=1;
					out<=238;
				end
				if(in == 631) begin
					state<=1;
					out<=239;
				end
				if(in == 632) begin
					state<=1;
					out<=240;
				end
				if(in == 633) begin
					state<=1;
					out<=241;
				end
				if(in == 634) begin
					state<=1;
					out<=242;
				end
				if(in == 635) begin
					state<=1;
					out<=243;
				end
				if(in == 636) begin
					state<=1;
					out<=244;
				end
				if(in == 637) begin
					state<=1;
					out<=245;
				end
				if(in == 638) begin
					state<=1;
					out<=246;
				end
				if(in == 639) begin
					state<=1;
					out<=247;
				end
				if(in == 640) begin
					state<=1;
					out<=248;
				end
				if(in == 641) begin
					state<=1;
					out<=249;
				end
				if(in == 642) begin
					state<=1;
					out<=250;
				end
				if(in == 643) begin
					state<=1;
					out<=251;
				end
				if(in == 644) begin
					state<=1;
					out<=252;
				end
				if(in == 645) begin
					state<=1;
					out<=253;
				end
				if(in == 646) begin
					state<=1;
					out<=254;
				end
				if(in == 647) begin
					state<=1;
					out<=255;
				end
				if(in == 648) begin
					state<=1;
					out<=0;
				end
				if(in == 649) begin
					state<=1;
					out<=1;
				end
				if(in == 650) begin
					state<=1;
					out<=2;
				end
				if(in == 651) begin
					state<=1;
					out<=3;
				end
				if(in == 652) begin
					state<=1;
					out<=4;
				end
				if(in == 653) begin
					state<=1;
					out<=5;
				end
				if(in == 654) begin
					state<=1;
					out<=6;
				end
				if(in == 655) begin
					state<=1;
					out<=7;
				end
				if(in == 656) begin
					state<=1;
					out<=8;
				end
				if(in == 657) begin
					state<=1;
					out<=9;
				end
				if(in == 658) begin
					state<=1;
					out<=10;
				end
				if(in == 659) begin
					state<=1;
					out<=11;
				end
				if(in == 660) begin
					state<=1;
					out<=12;
				end
				if(in == 661) begin
					state<=1;
					out<=13;
				end
				if(in == 662) begin
					state<=1;
					out<=14;
				end
				if(in == 663) begin
					state<=1;
					out<=15;
				end
				if(in == 664) begin
					state<=1;
					out<=16;
				end
				if(in == 665) begin
					state<=1;
					out<=17;
				end
				if(in == 666) begin
					state<=1;
					out<=18;
				end
				if(in == 667) begin
					state<=1;
					out<=19;
				end
				if(in == 668) begin
					state<=1;
					out<=20;
				end
				if(in == 669) begin
					state<=1;
					out<=21;
				end
				if(in == 670) begin
					state<=1;
					out<=22;
				end
				if(in == 671) begin
					state<=1;
					out<=23;
				end
				if(in == 672) begin
					state<=1;
					out<=24;
				end
				if(in == 673) begin
					state<=1;
					out<=25;
				end
				if(in == 674) begin
					state<=1;
					out<=26;
				end
				if(in == 675) begin
					state<=1;
					out<=27;
				end
				if(in == 676) begin
					state<=1;
					out<=28;
				end
				if(in == 677) begin
					state<=1;
					out<=29;
				end
				if(in == 678) begin
					state<=1;
					out<=30;
				end
				if(in == 679) begin
					state<=1;
					out<=31;
				end
				if(in == 680) begin
					state<=1;
					out<=32;
				end
				if(in == 681) begin
					state<=1;
					out<=33;
				end
				if(in == 682) begin
					state<=1;
					out<=34;
				end
				if(in == 683) begin
					state<=1;
					out<=35;
				end
				if(in == 684) begin
					state<=1;
					out<=36;
				end
				if(in == 685) begin
					state<=1;
					out<=37;
				end
				if(in == 686) begin
					state<=1;
					out<=38;
				end
				if(in == 687) begin
					state<=1;
					out<=39;
				end
				if(in == 688) begin
					state<=1;
					out<=40;
				end
				if(in == 689) begin
					state<=1;
					out<=41;
				end
				if(in == 690) begin
					state<=1;
					out<=42;
				end
				if(in == 691) begin
					state<=1;
					out<=43;
				end
				if(in == 692) begin
					state<=1;
					out<=44;
				end
				if(in == 693) begin
					state<=1;
					out<=45;
				end
				if(in == 694) begin
					state<=1;
					out<=46;
				end
				if(in == 695) begin
					state<=1;
					out<=47;
				end
				if(in == 696) begin
					state<=1;
					out<=48;
				end
				if(in == 697) begin
					state<=1;
					out<=49;
				end
				if(in == 698) begin
					state<=1;
					out<=50;
				end
				if(in == 699) begin
					state<=1;
					out<=51;
				end
				if(in == 700) begin
					state<=1;
					out<=52;
				end
				if(in == 701) begin
					state<=1;
					out<=53;
				end
				if(in == 702) begin
					state<=1;
					out<=54;
				end
				if(in == 703) begin
					state<=1;
					out<=55;
				end
				if(in == 704) begin
					state<=1;
					out<=56;
				end
				if(in == 705) begin
					state<=1;
					out<=57;
				end
				if(in == 706) begin
					state<=1;
					out<=58;
				end
				if(in == 707) begin
					state<=1;
					out<=59;
				end
				if(in == 708) begin
					state<=1;
					out<=60;
				end
				if(in == 709) begin
					state<=1;
					out<=61;
				end
				if(in == 710) begin
					state<=1;
					out<=62;
				end
				if(in == 711) begin
					state<=1;
					out<=63;
				end
				if(in == 712) begin
					state<=1;
					out<=64;
				end
				if(in == 713) begin
					state<=1;
					out<=65;
				end
				if(in == 714) begin
					state<=1;
					out<=66;
				end
				if(in == 715) begin
					state<=1;
					out<=67;
				end
				if(in == 716) begin
					state<=1;
					out<=68;
				end
				if(in == 717) begin
					state<=1;
					out<=69;
				end
				if(in == 718) begin
					state<=1;
					out<=70;
				end
				if(in == 719) begin
					state<=1;
					out<=71;
				end
				if(in == 720) begin
					state<=1;
					out<=72;
				end
				if(in == 721) begin
					state<=1;
					out<=73;
				end
				if(in == 722) begin
					state<=1;
					out<=74;
				end
				if(in == 723) begin
					state<=1;
					out<=75;
				end
				if(in == 724) begin
					state<=1;
					out<=76;
				end
				if(in == 725) begin
					state<=1;
					out<=77;
				end
				if(in == 726) begin
					state<=1;
					out<=78;
				end
				if(in == 727) begin
					state<=1;
					out<=79;
				end
				if(in == 728) begin
					state<=1;
					out<=80;
				end
				if(in == 729) begin
					state<=1;
					out<=81;
				end
				if(in == 730) begin
					state<=1;
					out<=82;
				end
				if(in == 731) begin
					state<=1;
					out<=83;
				end
				if(in == 732) begin
					state<=1;
					out<=84;
				end
				if(in == 733) begin
					state<=1;
					out<=85;
				end
				if(in == 734) begin
					state<=1;
					out<=86;
				end
				if(in == 735) begin
					state<=1;
					out<=87;
				end
				if(in == 736) begin
					state<=1;
					out<=88;
				end
				if(in == 737) begin
					state<=1;
					out<=89;
				end
				if(in == 738) begin
					state<=1;
					out<=90;
				end
				if(in == 739) begin
					state<=1;
					out<=91;
				end
				if(in == 740) begin
					state<=1;
					out<=92;
				end
				if(in == 741) begin
					state<=1;
					out<=93;
				end
				if(in == 742) begin
					state<=1;
					out<=94;
				end
				if(in == 743) begin
					state<=1;
					out<=95;
				end
				if(in == 744) begin
					state<=1;
					out<=96;
				end
				if(in == 745) begin
					state<=1;
					out<=97;
				end
				if(in == 746) begin
					state<=1;
					out<=98;
				end
				if(in == 747) begin
					state<=1;
					out<=99;
				end
				if(in == 748) begin
					state<=1;
					out<=100;
				end
				if(in == 749) begin
					state<=1;
					out<=101;
				end
				if(in == 750) begin
					state<=1;
					out<=102;
				end
				if(in == 751) begin
					state<=1;
					out<=103;
				end
				if(in == 752) begin
					state<=1;
					out<=104;
				end
				if(in == 753) begin
					state<=1;
					out<=105;
				end
				if(in == 754) begin
					state<=1;
					out<=106;
				end
				if(in == 755) begin
					state<=1;
					out<=107;
				end
				if(in == 756) begin
					state<=1;
					out<=108;
				end
				if(in == 757) begin
					state<=1;
					out<=109;
				end
				if(in == 758) begin
					state<=1;
					out<=110;
				end
				if(in == 759) begin
					state<=1;
					out<=111;
				end
				if(in == 760) begin
					state<=1;
					out<=112;
				end
				if(in == 761) begin
					state<=1;
					out<=113;
				end
				if(in == 762) begin
					state<=1;
					out<=114;
				end
				if(in == 763) begin
					state<=1;
					out<=115;
				end
				if(in == 764) begin
					state<=1;
					out<=116;
				end
				if(in == 765) begin
					state<=1;
					out<=117;
				end
				if(in == 766) begin
					state<=1;
					out<=118;
				end
				if(in == 767) begin
					state<=1;
					out<=119;
				end
				if(in == 768) begin
					state<=1;
					out<=120;
				end
				if(in == 769) begin
					state<=1;
					out<=121;
				end
				if(in == 770) begin
					state<=1;
					out<=122;
				end
				if(in == 771) begin
					state<=1;
					out<=123;
				end
				if(in == 772) begin
					state<=1;
					out<=124;
				end
				if(in == 773) begin
					state<=1;
					out<=125;
				end
				if(in == 774) begin
					state<=1;
					out<=126;
				end
				if(in == 775) begin
					state<=1;
					out<=127;
				end
				if(in == 776) begin
					state<=1;
					out<=128;
				end
				if(in == 777) begin
					state<=1;
					out<=129;
				end
				if(in == 778) begin
					state<=1;
					out<=130;
				end
				if(in == 779) begin
					state<=1;
					out<=131;
				end
				if(in == 780) begin
					state<=1;
					out<=132;
				end
				if(in == 781) begin
					state<=1;
					out<=133;
				end
				if(in == 782) begin
					state<=1;
					out<=134;
				end
				if(in == 783) begin
					state<=1;
					out<=135;
				end
				if(in == 784) begin
					state<=1;
					out<=136;
				end
				if(in == 785) begin
					state<=1;
					out<=137;
				end
				if(in == 786) begin
					state<=1;
					out<=138;
				end
				if(in == 787) begin
					state<=1;
					out<=139;
				end
				if(in == 788) begin
					state<=1;
					out<=140;
				end
				if(in == 789) begin
					state<=1;
					out<=141;
				end
				if(in == 790) begin
					state<=1;
					out<=142;
				end
				if(in == 791) begin
					state<=1;
					out<=143;
				end
				if(in == 792) begin
					state<=1;
					out<=144;
				end
				if(in == 793) begin
					state<=1;
					out<=145;
				end
				if(in == 794) begin
					state<=1;
					out<=146;
				end
				if(in == 795) begin
					state<=1;
					out<=147;
				end
				if(in == 796) begin
					state<=1;
					out<=148;
				end
				if(in == 797) begin
					state<=1;
					out<=149;
				end
				if(in == 798) begin
					state<=1;
					out<=150;
				end
				if(in == 799) begin
					state<=1;
					out<=151;
				end
				if(in == 800) begin
					state<=1;
					out<=152;
				end
				if(in == 801) begin
					state<=1;
					out<=153;
				end
				if(in == 802) begin
					state<=1;
					out<=154;
				end
				if(in == 803) begin
					state<=1;
					out<=155;
				end
				if(in == 804) begin
					state<=1;
					out<=156;
				end
				if(in == 805) begin
					state<=1;
					out<=157;
				end
				if(in == 806) begin
					state<=1;
					out<=158;
				end
				if(in == 807) begin
					state<=1;
					out<=159;
				end
				if(in == 808) begin
					state<=1;
					out<=160;
				end
				if(in == 809) begin
					state<=1;
					out<=161;
				end
				if(in == 810) begin
					state<=1;
					out<=162;
				end
				if(in == 811) begin
					state<=1;
					out<=163;
				end
				if(in == 812) begin
					state<=1;
					out<=164;
				end
				if(in == 813) begin
					state<=1;
					out<=165;
				end
				if(in == 814) begin
					state<=1;
					out<=166;
				end
				if(in == 815) begin
					state<=1;
					out<=167;
				end
				if(in == 816) begin
					state<=1;
					out<=168;
				end
				if(in == 817) begin
					state<=1;
					out<=169;
				end
				if(in == 818) begin
					state<=1;
					out<=170;
				end
				if(in == 819) begin
					state<=1;
					out<=171;
				end
				if(in == 820) begin
					state<=1;
					out<=172;
				end
				if(in == 821) begin
					state<=1;
					out<=173;
				end
				if(in == 822) begin
					state<=1;
					out<=174;
				end
				if(in == 823) begin
					state<=1;
					out<=175;
				end
				if(in == 824) begin
					state<=1;
					out<=176;
				end
				if(in == 825) begin
					state<=1;
					out<=177;
				end
				if(in == 826) begin
					state<=1;
					out<=178;
				end
				if(in == 827) begin
					state<=1;
					out<=179;
				end
				if(in == 828) begin
					state<=1;
					out<=180;
				end
				if(in == 829) begin
					state<=1;
					out<=181;
				end
				if(in == 830) begin
					state<=1;
					out<=182;
				end
				if(in == 831) begin
					state<=1;
					out<=183;
				end
				if(in == 832) begin
					state<=1;
					out<=184;
				end
				if(in == 833) begin
					state<=1;
					out<=185;
				end
				if(in == 834) begin
					state<=1;
					out<=186;
				end
				if(in == 835) begin
					state<=1;
					out<=187;
				end
				if(in == 836) begin
					state<=1;
					out<=188;
				end
				if(in == 837) begin
					state<=1;
					out<=189;
				end
				if(in == 838) begin
					state<=1;
					out<=190;
				end
				if(in == 839) begin
					state<=1;
					out<=191;
				end
				if(in == 840) begin
					state<=1;
					out<=192;
				end
				if(in == 841) begin
					state<=1;
					out<=193;
				end
				if(in == 842) begin
					state<=1;
					out<=194;
				end
				if(in == 843) begin
					state<=1;
					out<=195;
				end
				if(in == 844) begin
					state<=1;
					out<=196;
				end
				if(in == 845) begin
					state<=1;
					out<=197;
				end
				if(in == 846) begin
					state<=1;
					out<=198;
				end
				if(in == 847) begin
					state<=1;
					out<=199;
				end
				if(in == 848) begin
					state<=1;
					out<=200;
				end
				if(in == 849) begin
					state<=1;
					out<=201;
				end
				if(in == 850) begin
					state<=1;
					out<=202;
				end
				if(in == 851) begin
					state<=1;
					out<=203;
				end
				if(in == 852) begin
					state<=1;
					out<=204;
				end
				if(in == 853) begin
					state<=1;
					out<=205;
				end
				if(in == 854) begin
					state<=1;
					out<=206;
				end
				if(in == 855) begin
					state<=1;
					out<=207;
				end
				if(in == 856) begin
					state<=1;
					out<=208;
				end
				if(in == 857) begin
					state<=1;
					out<=209;
				end
				if(in == 858) begin
					state<=1;
					out<=210;
				end
				if(in == 859) begin
					state<=1;
					out<=211;
				end
				if(in == 860) begin
					state<=1;
					out<=212;
				end
				if(in == 861) begin
					state<=1;
					out<=213;
				end
				if(in == 862) begin
					state<=1;
					out<=214;
				end
				if(in == 863) begin
					state<=1;
					out<=215;
				end
				if(in == 864) begin
					state<=1;
					out<=216;
				end
				if(in == 865) begin
					state<=1;
					out<=217;
				end
				if(in == 866) begin
					state<=1;
					out<=218;
				end
				if(in == 867) begin
					state<=1;
					out<=219;
				end
				if(in == 868) begin
					state<=1;
					out<=220;
				end
				if(in == 869) begin
					state<=1;
					out<=221;
				end
				if(in == 870) begin
					state<=1;
					out<=222;
				end
				if(in == 871) begin
					state<=1;
					out<=223;
				end
				if(in == 872) begin
					state<=1;
					out<=224;
				end
				if(in == 873) begin
					state<=1;
					out<=225;
				end
				if(in == 874) begin
					state<=1;
					out<=226;
				end
				if(in == 875) begin
					state<=1;
					out<=227;
				end
				if(in == 876) begin
					state<=1;
					out<=228;
				end
				if(in == 877) begin
					state<=1;
					out<=229;
				end
				if(in == 878) begin
					state<=1;
					out<=230;
				end
				if(in == 879) begin
					state<=1;
					out<=231;
				end
				if(in == 880) begin
					state<=1;
					out<=232;
				end
				if(in == 881) begin
					state<=1;
					out<=233;
				end
				if(in == 882) begin
					state<=1;
					out<=234;
				end
				if(in == 883) begin
					state<=1;
					out<=235;
				end
				if(in == 884) begin
					state<=1;
					out<=236;
				end
				if(in == 885) begin
					state<=1;
					out<=237;
				end
				if(in == 886) begin
					state<=1;
					out<=238;
				end
				if(in == 887) begin
					state<=1;
					out<=239;
				end
				if(in == 888) begin
					state<=1;
					out<=240;
				end
				if(in == 889) begin
					state<=1;
					out<=241;
				end
				if(in == 890) begin
					state<=1;
					out<=242;
				end
				if(in == 891) begin
					state<=1;
					out<=243;
				end
				if(in == 892) begin
					state<=1;
					out<=244;
				end
				if(in == 893) begin
					state<=1;
					out<=245;
				end
				if(in == 894) begin
					state<=1;
					out<=246;
				end
				if(in == 895) begin
					state<=1;
					out<=247;
				end
				if(in == 896) begin
					state<=1;
					out<=248;
				end
				if(in == 897) begin
					state<=1;
					out<=249;
				end
				if(in == 898) begin
					state<=1;
					out<=250;
				end
				if(in == 899) begin
					state<=1;
					out<=251;
				end
				if(in == 900) begin
					state<=1;
					out<=252;
				end
				if(in == 901) begin
					state<=1;
					out<=253;
				end
				if(in == 902) begin
					state<=1;
					out<=254;
				end
				if(in == 903) begin
					state<=1;
					out<=255;
				end
				if(in == 904) begin
					state<=1;
					out<=0;
				end
				if(in == 905) begin
					state<=1;
					out<=1;
				end
				if(in == 906) begin
					state<=1;
					out<=2;
				end
				if(in == 907) begin
					state<=1;
					out<=3;
				end
				if(in == 908) begin
					state<=1;
					out<=4;
				end
				if(in == 909) begin
					state<=1;
					out<=5;
				end
				if(in == 910) begin
					state<=1;
					out<=6;
				end
				if(in == 911) begin
					state<=1;
					out<=7;
				end
				if(in == 912) begin
					state<=1;
					out<=8;
				end
				if(in == 913) begin
					state<=1;
					out<=9;
				end
				if(in == 914) begin
					state<=1;
					out<=10;
				end
				if(in == 915) begin
					state<=1;
					out<=11;
				end
				if(in == 916) begin
					state<=1;
					out<=12;
				end
				if(in == 917) begin
					state<=1;
					out<=13;
				end
				if(in == 918) begin
					state<=1;
					out<=14;
				end
				if(in == 919) begin
					state<=1;
					out<=15;
				end
				if(in == 920) begin
					state<=1;
					out<=16;
				end
				if(in == 921) begin
					state<=1;
					out<=17;
				end
				if(in == 922) begin
					state<=1;
					out<=18;
				end
				if(in == 923) begin
					state<=1;
					out<=19;
				end
				if(in == 924) begin
					state<=1;
					out<=20;
				end
				if(in == 925) begin
					state<=1;
					out<=21;
				end
				if(in == 926) begin
					state<=1;
					out<=22;
				end
				if(in == 927) begin
					state<=1;
					out<=23;
				end
				if(in == 928) begin
					state<=1;
					out<=24;
				end
			end
		endcase
	end
endmodule