module s27();