module s382(input clk,input[2:0] in, output [7:0] out);
	reg[12:0] state;
	always @(posedge clk) begin
		out<=0;
		case (state)
			0: begin
				if(in == 0) begin
					state<=800;
					out<=0;
				end
				if(in == 1) begin
					state<=1231;
					out<=1;
				end
				if(in == 2) begin
					state<=2621;
					out<=2;
				end
				if(in == 3) begin
					state<=5129;
					out<=3;
				end
				if(in == 4) begin
					state<=6510;
					out<=4;
				end
			end
			1: begin
				if(in == 0) begin
					state<=2;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=3900;
					out<=7;
				end
				if(in == 3) begin
					state<=2000;
					out<=8;
				end
				if(in == 4) begin
					state<=5889;
					out<=9;
				end
			end
			2: begin
				if(in == 0) begin
					state<=3;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=3901;
					out<=12;
				end
				if(in == 3) begin
					state<=2001;
					out<=13;
				end
				if(in == 4) begin
					state<=5890;
					out<=14;
				end
			end
			3: begin
				if(in == 0) begin
					state<=4;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=3902;
					out<=17;
				end
				if(in == 3) begin
					state<=2002;
					out<=18;
				end
				if(in == 4) begin
					state<=5891;
					out<=19;
				end
			end
			4: begin
				if(in == 0) begin
					state<=5;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=3903;
					out<=22;
				end
				if(in == 3) begin
					state<=2003;
					out<=23;
				end
				if(in == 4) begin
					state<=5892;
					out<=24;
				end
			end
			5: begin
				if(in == 0) begin
					state<=6;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=3904;
					out<=27;
				end
				if(in == 3) begin
					state<=2004;
					out<=28;
				end
				if(in == 4) begin
					state<=5893;
					out<=29;
				end
			end
			6: begin
				if(in == 0) begin
					state<=7;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=3905;
					out<=32;
				end
				if(in == 3) begin
					state<=2005;
					out<=33;
				end
				if(in == 4) begin
					state<=5894;
					out<=34;
				end
			end
			7: begin
				if(in == 0) begin
					state<=8;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=3906;
					out<=37;
				end
				if(in == 3) begin
					state<=2006;
					out<=38;
				end
				if(in == 4) begin
					state<=5895;
					out<=39;
				end
			end
			8: begin
				if(in == 0) begin
					state<=9;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=3907;
					out<=42;
				end
				if(in == 3) begin
					state<=2007;
					out<=43;
				end
				if(in == 4) begin
					state<=5896;
					out<=44;
				end
			end
			9: begin
				if(in == 0) begin
					state<=10;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=3908;
					out<=47;
				end
				if(in == 3) begin
					state<=2008;
					out<=48;
				end
				if(in == 4) begin
					state<=5897;
					out<=49;
				end
			end
			10: begin
				if(in == 0) begin
					state<=11;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=3909;
					out<=52;
				end
				if(in == 3) begin
					state<=2009;
					out<=53;
				end
				if(in == 4) begin
					state<=5898;
					out<=54;
				end
			end
			11: begin
				if(in == 0) begin
					state<=12;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=3910;
					out<=57;
				end
				if(in == 3) begin
					state<=2010;
					out<=58;
				end
				if(in == 4) begin
					state<=5899;
					out<=59;
				end
			end
			12: begin
				if(in == 0) begin
					state<=13;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=3911;
					out<=62;
				end
				if(in == 3) begin
					state<=2011;
					out<=63;
				end
				if(in == 4) begin
					state<=5900;
					out<=64;
				end
			end
			13: begin
				if(in == 0) begin
					state<=14;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=3912;
					out<=67;
				end
				if(in == 3) begin
					state<=2012;
					out<=68;
				end
				if(in == 4) begin
					state<=5901;
					out<=69;
				end
			end
			14: begin
				if(in == 0) begin
					state<=15;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=3913;
					out<=72;
				end
				if(in == 3) begin
					state<=2013;
					out<=73;
				end
				if(in == 4) begin
					state<=5902;
					out<=74;
				end
			end
			15: begin
				if(in == 0) begin
					state<=16;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=3914;
					out<=77;
				end
				if(in == 3) begin
					state<=2014;
					out<=78;
				end
				if(in == 4) begin
					state<=5903;
					out<=79;
				end
			end
			16: begin
				if(in == 0) begin
					state<=17;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=3915;
					out<=82;
				end
				if(in == 3) begin
					state<=2015;
					out<=83;
				end
				if(in == 4) begin
					state<=5904;
					out<=84;
				end
			end
			17: begin
				if(in == 0) begin
					state<=18;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=3916;
					out<=87;
				end
				if(in == 3) begin
					state<=2016;
					out<=88;
				end
				if(in == 4) begin
					state<=5905;
					out<=89;
				end
			end
			18: begin
				if(in == 0) begin
					state<=19;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=3917;
					out<=92;
				end
				if(in == 3) begin
					state<=2017;
					out<=93;
				end
				if(in == 4) begin
					state<=5906;
					out<=94;
				end
			end
			19: begin
				if(in == 0) begin
					state<=20;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=3918;
					out<=97;
				end
				if(in == 3) begin
					state<=2018;
					out<=98;
				end
				if(in == 4) begin
					state<=5907;
					out<=99;
				end
			end
			20: begin
				if(in == 0) begin
					state<=21;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=3919;
					out<=102;
				end
				if(in == 3) begin
					state<=2019;
					out<=103;
				end
				if(in == 4) begin
					state<=5908;
					out<=104;
				end
			end
			21: begin
				if(in == 0) begin
					state<=22;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=3920;
					out<=107;
				end
				if(in == 3) begin
					state<=2020;
					out<=108;
				end
				if(in == 4) begin
					state<=5909;
					out<=109;
				end
			end
			22: begin
				if(in == 0) begin
					state<=23;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=3921;
					out<=112;
				end
				if(in == 3) begin
					state<=2021;
					out<=113;
				end
				if(in == 4) begin
					state<=5910;
					out<=114;
				end
			end
			23: begin
				if(in == 0) begin
					state<=24;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=3922;
					out<=117;
				end
				if(in == 3) begin
					state<=2022;
					out<=118;
				end
				if(in == 4) begin
					state<=5911;
					out<=119;
				end
			end
			24: begin
				if(in == 0) begin
					state<=25;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=3923;
					out<=122;
				end
				if(in == 3) begin
					state<=2023;
					out<=123;
				end
				if(in == 4) begin
					state<=5912;
					out<=124;
				end
			end
			25: begin
				if(in == 0) begin
					state<=26;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=3924;
					out<=127;
				end
				if(in == 3) begin
					state<=2024;
					out<=128;
				end
				if(in == 4) begin
					state<=5913;
					out<=129;
				end
			end
			26: begin
				if(in == 0) begin
					state<=27;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=3925;
					out<=132;
				end
				if(in == 3) begin
					state<=2025;
					out<=133;
				end
				if(in == 4) begin
					state<=5914;
					out<=134;
				end
			end
			27: begin
				if(in == 0) begin
					state<=28;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=3926;
					out<=137;
				end
				if(in == 3) begin
					state<=2026;
					out<=138;
				end
				if(in == 4) begin
					state<=5915;
					out<=139;
				end
			end
			28: begin
				if(in == 0) begin
					state<=29;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=3927;
					out<=142;
				end
				if(in == 3) begin
					state<=2027;
					out<=143;
				end
				if(in == 4) begin
					state<=5916;
					out<=144;
				end
			end
			29: begin
				if(in == 0) begin
					state<=30;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=3928;
					out<=147;
				end
				if(in == 3) begin
					state<=2028;
					out<=148;
				end
				if(in == 4) begin
					state<=5917;
					out<=149;
				end
			end
			30: begin
				if(in == 0) begin
					state<=31;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=3929;
					out<=152;
				end
				if(in == 3) begin
					state<=2029;
					out<=153;
				end
				if(in == 4) begin
					state<=5918;
					out<=154;
				end
			end
			31: begin
				if(in == 0) begin
					state<=32;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=3930;
					out<=157;
				end
				if(in == 3) begin
					state<=2030;
					out<=158;
				end
				if(in == 4) begin
					state<=5919;
					out<=159;
				end
			end
			32: begin
				if(in == 0) begin
					state<=33;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=3931;
					out<=162;
				end
				if(in == 3) begin
					state<=2031;
					out<=163;
				end
				if(in == 4) begin
					state<=5920;
					out<=164;
				end
			end
			33: begin
				if(in == 0) begin
					state<=34;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=3932;
					out<=167;
				end
				if(in == 3) begin
					state<=2032;
					out<=168;
				end
				if(in == 4) begin
					state<=5921;
					out<=169;
				end
			end
			34: begin
				if(in == 0) begin
					state<=35;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=3933;
					out<=172;
				end
				if(in == 3) begin
					state<=2033;
					out<=173;
				end
				if(in == 4) begin
					state<=5922;
					out<=174;
				end
			end
			35: begin
				if(in == 0) begin
					state<=36;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=3934;
					out<=177;
				end
				if(in == 3) begin
					state<=2034;
					out<=178;
				end
				if(in == 4) begin
					state<=5923;
					out<=179;
				end
			end
			36: begin
				if(in == 0) begin
					state<=37;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=3935;
					out<=182;
				end
				if(in == 3) begin
					state<=2035;
					out<=183;
				end
				if(in == 4) begin
					state<=5924;
					out<=184;
				end
			end
			37: begin
				if(in == 0) begin
					state<=38;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=3936;
					out<=187;
				end
				if(in == 3) begin
					state<=2036;
					out<=188;
				end
				if(in == 4) begin
					state<=5925;
					out<=189;
				end
			end
			38: begin
				if(in == 0) begin
					state<=39;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=3937;
					out<=192;
				end
				if(in == 3) begin
					state<=2037;
					out<=193;
				end
				if(in == 4) begin
					state<=5926;
					out<=194;
				end
			end
			39: begin
				if(in == 0) begin
					state<=40;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=3938;
					out<=197;
				end
				if(in == 3) begin
					state<=2038;
					out<=198;
				end
				if(in == 4) begin
					state<=5927;
					out<=199;
				end
			end
			40: begin
				if(in == 0) begin
					state<=41;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=3939;
					out<=202;
				end
				if(in == 3) begin
					state<=2039;
					out<=203;
				end
				if(in == 4) begin
					state<=5928;
					out<=204;
				end
			end
			41: begin
				if(in == 0) begin
					state<=42;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=3940;
					out<=207;
				end
				if(in == 3) begin
					state<=2040;
					out<=208;
				end
				if(in == 4) begin
					state<=5929;
					out<=209;
				end
			end
			42: begin
				if(in == 0) begin
					state<=43;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=3941;
					out<=212;
				end
				if(in == 3) begin
					state<=2041;
					out<=213;
				end
				if(in == 4) begin
					state<=5930;
					out<=214;
				end
			end
			43: begin
				if(in == 0) begin
					state<=44;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=3942;
					out<=217;
				end
				if(in == 3) begin
					state<=2042;
					out<=218;
				end
				if(in == 4) begin
					state<=5931;
					out<=219;
				end
			end
			44: begin
				if(in == 0) begin
					state<=45;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=3943;
					out<=222;
				end
				if(in == 3) begin
					state<=2043;
					out<=223;
				end
				if(in == 4) begin
					state<=5932;
					out<=224;
				end
			end
			45: begin
				if(in == 0) begin
					state<=46;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=3944;
					out<=227;
				end
				if(in == 3) begin
					state<=2044;
					out<=228;
				end
				if(in == 4) begin
					state<=5933;
					out<=229;
				end
			end
			46: begin
				if(in == 0) begin
					state<=47;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=3945;
					out<=232;
				end
				if(in == 3) begin
					state<=2045;
					out<=233;
				end
				if(in == 4) begin
					state<=5934;
					out<=234;
				end
			end
			47: begin
				if(in == 0) begin
					state<=48;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=3946;
					out<=237;
				end
				if(in == 3) begin
					state<=2046;
					out<=238;
				end
				if(in == 4) begin
					state<=5935;
					out<=239;
				end
			end
			48: begin
				if(in == 0) begin
					state<=49;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=3947;
					out<=242;
				end
				if(in == 3) begin
					state<=2047;
					out<=243;
				end
				if(in == 4) begin
					state<=5936;
					out<=244;
				end
			end
			49: begin
				if(in == 0) begin
					state<=50;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=3948;
					out<=247;
				end
				if(in == 3) begin
					state<=2048;
					out<=248;
				end
				if(in == 4) begin
					state<=5937;
					out<=249;
				end
			end
			50: begin
				if(in == 0) begin
					state<=1329;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=5218;
					out<=252;
				end
				if(in == 3) begin
					state<=3261;
					out<=253;
				end
				if(in == 4) begin
					state<=7150;
					out<=254;
				end
			end
			51: begin
				if(in == 0) begin
					state<=52;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=3950;
					out<=1;
				end
				if(in == 3) begin
					state<=2050;
					out<=2;
				end
				if(in == 4) begin
					state<=5939;
					out<=3;
				end
			end
			52: begin
				if(in == 0) begin
					state<=53;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=3951;
					out<=6;
				end
				if(in == 3) begin
					state<=2051;
					out<=7;
				end
				if(in == 4) begin
					state<=5940;
					out<=8;
				end
			end
			53: begin
				if(in == 0) begin
					state<=54;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=3952;
					out<=11;
				end
				if(in == 3) begin
					state<=2052;
					out<=12;
				end
				if(in == 4) begin
					state<=5941;
					out<=13;
				end
			end
			54: begin
				if(in == 0) begin
					state<=55;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=3953;
					out<=16;
				end
				if(in == 3) begin
					state<=2053;
					out<=17;
				end
				if(in == 4) begin
					state<=5942;
					out<=18;
				end
			end
			55: begin
				if(in == 0) begin
					state<=56;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=3954;
					out<=21;
				end
				if(in == 3) begin
					state<=2054;
					out<=22;
				end
				if(in == 4) begin
					state<=5943;
					out<=23;
				end
			end
			56: begin
				if(in == 0) begin
					state<=57;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=3955;
					out<=26;
				end
				if(in == 3) begin
					state<=2055;
					out<=27;
				end
				if(in == 4) begin
					state<=5944;
					out<=28;
				end
			end
			57: begin
				if(in == 0) begin
					state<=58;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=3956;
					out<=31;
				end
				if(in == 3) begin
					state<=2056;
					out<=32;
				end
				if(in == 4) begin
					state<=5945;
					out<=33;
				end
			end
			58: begin
				if(in == 0) begin
					state<=59;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=3957;
					out<=36;
				end
				if(in == 3) begin
					state<=2057;
					out<=37;
				end
				if(in == 4) begin
					state<=5946;
					out<=38;
				end
			end
			59: begin
				if(in == 0) begin
					state<=60;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=3958;
					out<=41;
				end
				if(in == 3) begin
					state<=2058;
					out<=42;
				end
				if(in == 4) begin
					state<=5947;
					out<=43;
				end
			end
			60: begin
				if(in == 0) begin
					state<=61;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=3959;
					out<=46;
				end
				if(in == 3) begin
					state<=2059;
					out<=47;
				end
				if(in == 4) begin
					state<=5948;
					out<=48;
				end
			end
			61: begin
				if(in == 0) begin
					state<=62;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=3960;
					out<=51;
				end
				if(in == 3) begin
					state<=2060;
					out<=52;
				end
				if(in == 4) begin
					state<=5949;
					out<=53;
				end
			end
			62: begin
				if(in == 0) begin
					state<=63;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=3961;
					out<=56;
				end
				if(in == 3) begin
					state<=2061;
					out<=57;
				end
				if(in == 4) begin
					state<=5950;
					out<=58;
				end
			end
			63: begin
				if(in == 0) begin
					state<=64;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=3962;
					out<=61;
				end
				if(in == 3) begin
					state<=2062;
					out<=62;
				end
				if(in == 4) begin
					state<=5951;
					out<=63;
				end
			end
			64: begin
				if(in == 0) begin
					state<=65;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=3963;
					out<=66;
				end
				if(in == 3) begin
					state<=2063;
					out<=67;
				end
				if(in == 4) begin
					state<=5952;
					out<=68;
				end
			end
			65: begin
				if(in == 0) begin
					state<=66;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=3964;
					out<=71;
				end
				if(in == 3) begin
					state<=2064;
					out<=72;
				end
				if(in == 4) begin
					state<=5953;
					out<=73;
				end
			end
			66: begin
				if(in == 0) begin
					state<=67;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=3965;
					out<=76;
				end
				if(in == 3) begin
					state<=2065;
					out<=77;
				end
				if(in == 4) begin
					state<=5954;
					out<=78;
				end
			end
			67: begin
				if(in == 0) begin
					state<=68;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=3966;
					out<=81;
				end
				if(in == 3) begin
					state<=2066;
					out<=82;
				end
				if(in == 4) begin
					state<=5955;
					out<=83;
				end
			end
			68: begin
				if(in == 0) begin
					state<=69;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=3967;
					out<=86;
				end
				if(in == 3) begin
					state<=2067;
					out<=87;
				end
				if(in == 4) begin
					state<=5956;
					out<=88;
				end
			end
			69: begin
				if(in == 0) begin
					state<=70;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=3968;
					out<=91;
				end
				if(in == 3) begin
					state<=2068;
					out<=92;
				end
				if(in == 4) begin
					state<=5957;
					out<=93;
				end
			end
			70: begin
				if(in == 0) begin
					state<=71;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=3969;
					out<=96;
				end
				if(in == 3) begin
					state<=2069;
					out<=97;
				end
				if(in == 4) begin
					state<=5958;
					out<=98;
				end
			end
			71: begin
				if(in == 0) begin
					state<=72;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=3970;
					out<=101;
				end
				if(in == 3) begin
					state<=2070;
					out<=102;
				end
				if(in == 4) begin
					state<=5959;
					out<=103;
				end
			end
			72: begin
				if(in == 0) begin
					state<=73;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=3971;
					out<=106;
				end
				if(in == 3) begin
					state<=2071;
					out<=107;
				end
				if(in == 4) begin
					state<=5960;
					out<=108;
				end
			end
			73: begin
				if(in == 0) begin
					state<=74;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=3972;
					out<=111;
				end
				if(in == 3) begin
					state<=2072;
					out<=112;
				end
				if(in == 4) begin
					state<=5961;
					out<=113;
				end
			end
			74: begin
				if(in == 0) begin
					state<=75;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=3973;
					out<=116;
				end
				if(in == 3) begin
					state<=2073;
					out<=117;
				end
				if(in == 4) begin
					state<=5962;
					out<=118;
				end
			end
			75: begin
				if(in == 0) begin
					state<=76;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=3974;
					out<=121;
				end
				if(in == 3) begin
					state<=2074;
					out<=122;
				end
				if(in == 4) begin
					state<=5963;
					out<=123;
				end
			end
			76: begin
				if(in == 0) begin
					state<=77;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=3975;
					out<=126;
				end
				if(in == 3) begin
					state<=2075;
					out<=127;
				end
				if(in == 4) begin
					state<=5964;
					out<=128;
				end
			end
			77: begin
				if(in == 0) begin
					state<=78;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=3976;
					out<=131;
				end
				if(in == 3) begin
					state<=2076;
					out<=132;
				end
				if(in == 4) begin
					state<=5965;
					out<=133;
				end
			end
			78: begin
				if(in == 0) begin
					state<=79;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=3977;
					out<=136;
				end
				if(in == 3) begin
					state<=2077;
					out<=137;
				end
				if(in == 4) begin
					state<=5966;
					out<=138;
				end
			end
			79: begin
				if(in == 0) begin
					state<=80;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=3978;
					out<=141;
				end
				if(in == 3) begin
					state<=2078;
					out<=142;
				end
				if(in == 4) begin
					state<=5967;
					out<=143;
				end
			end
			80: begin
				if(in == 0) begin
					state<=81;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=3979;
					out<=146;
				end
				if(in == 3) begin
					state<=2079;
					out<=147;
				end
				if(in == 4) begin
					state<=5968;
					out<=148;
				end
			end
			81: begin
				if(in == 0) begin
					state<=82;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=3980;
					out<=151;
				end
				if(in == 3) begin
					state<=2080;
					out<=152;
				end
				if(in == 4) begin
					state<=5969;
					out<=153;
				end
			end
			82: begin
				if(in == 0) begin
					state<=83;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=3981;
					out<=156;
				end
				if(in == 3) begin
					state<=2081;
					out<=157;
				end
				if(in == 4) begin
					state<=5970;
					out<=158;
				end
			end
			83: begin
				if(in == 0) begin
					state<=84;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=3982;
					out<=161;
				end
				if(in == 3) begin
					state<=2082;
					out<=162;
				end
				if(in == 4) begin
					state<=5971;
					out<=163;
				end
			end
			84: begin
				if(in == 0) begin
					state<=85;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=3983;
					out<=166;
				end
				if(in == 3) begin
					state<=2083;
					out<=167;
				end
				if(in == 4) begin
					state<=5972;
					out<=168;
				end
			end
			85: begin
				if(in == 0) begin
					state<=86;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=3984;
					out<=171;
				end
				if(in == 3) begin
					state<=2084;
					out<=172;
				end
				if(in == 4) begin
					state<=5973;
					out<=173;
				end
			end
			86: begin
				if(in == 0) begin
					state<=87;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=3985;
					out<=176;
				end
				if(in == 3) begin
					state<=2085;
					out<=177;
				end
				if(in == 4) begin
					state<=5974;
					out<=178;
				end
			end
			87: begin
				if(in == 0) begin
					state<=88;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=3986;
					out<=181;
				end
				if(in == 3) begin
					state<=2086;
					out<=182;
				end
				if(in == 4) begin
					state<=5975;
					out<=183;
				end
			end
			88: begin
				if(in == 0) begin
					state<=89;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=3987;
					out<=186;
				end
				if(in == 3) begin
					state<=2087;
					out<=187;
				end
				if(in == 4) begin
					state<=5976;
					out<=188;
				end
			end
			89: begin
				if(in == 0) begin
					state<=90;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=3988;
					out<=191;
				end
				if(in == 3) begin
					state<=2088;
					out<=192;
				end
				if(in == 4) begin
					state<=5977;
					out<=193;
				end
			end
			90: begin
				if(in == 0) begin
					state<=91;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=3989;
					out<=196;
				end
				if(in == 3) begin
					state<=2089;
					out<=197;
				end
				if(in == 4) begin
					state<=5978;
					out<=198;
				end
			end
			91: begin
				if(in == 0) begin
					state<=92;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=3990;
					out<=201;
				end
				if(in == 3) begin
					state<=2090;
					out<=202;
				end
				if(in == 4) begin
					state<=5979;
					out<=203;
				end
			end
			92: begin
				if(in == 0) begin
					state<=93;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=3991;
					out<=206;
				end
				if(in == 3) begin
					state<=2091;
					out<=207;
				end
				if(in == 4) begin
					state<=5980;
					out<=208;
				end
			end
			93: begin
				if(in == 0) begin
					state<=94;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=3992;
					out<=211;
				end
				if(in == 3) begin
					state<=2092;
					out<=212;
				end
				if(in == 4) begin
					state<=5981;
					out<=213;
				end
			end
			94: begin
				if(in == 0) begin
					state<=95;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=3993;
					out<=216;
				end
				if(in == 3) begin
					state<=2093;
					out<=217;
				end
				if(in == 4) begin
					state<=5982;
					out<=218;
				end
			end
			95: begin
				if(in == 0) begin
					state<=96;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=3994;
					out<=221;
				end
				if(in == 3) begin
					state<=2094;
					out<=222;
				end
				if(in == 4) begin
					state<=5983;
					out<=223;
				end
			end
			96: begin
				if(in == 0) begin
					state<=97;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=3995;
					out<=226;
				end
				if(in == 3) begin
					state<=2095;
					out<=227;
				end
				if(in == 4) begin
					state<=5984;
					out<=228;
				end
			end
			97: begin
				if(in == 0) begin
					state<=98;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=3996;
					out<=231;
				end
				if(in == 3) begin
					state<=2096;
					out<=232;
				end
				if(in == 4) begin
					state<=5985;
					out<=233;
				end
			end
			98: begin
				if(in == 0) begin
					state<=99;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=3997;
					out<=236;
				end
				if(in == 3) begin
					state<=2097;
					out<=237;
				end
				if(in == 4) begin
					state<=5986;
					out<=238;
				end
			end
			99: begin
				if(in == 0) begin
					state<=100;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=3998;
					out<=241;
				end
				if(in == 3) begin
					state<=2098;
					out<=242;
				end
				if(in == 4) begin
					state<=5987;
					out<=243;
				end
			end
			100: begin
				if(in == 0) begin
					state<=101;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=3999;
					out<=246;
				end
				if(in == 3) begin
					state<=2099;
					out<=247;
				end
				if(in == 4) begin
					state<=5988;
					out<=248;
				end
			end
			101: begin
				if(in == 0) begin
					state<=102;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=4000;
					out<=251;
				end
				if(in == 3) begin
					state<=2100;
					out<=252;
				end
				if(in == 4) begin
					state<=5989;
					out<=253;
				end
			end
			102: begin
				if(in == 0) begin
					state<=103;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=4001;
					out<=0;
				end
				if(in == 3) begin
					state<=2101;
					out<=1;
				end
				if(in == 4) begin
					state<=5990;
					out<=2;
				end
			end
			103: begin
				if(in == 0) begin
					state<=104;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=4002;
					out<=5;
				end
				if(in == 3) begin
					state<=2102;
					out<=6;
				end
				if(in == 4) begin
					state<=5991;
					out<=7;
				end
			end
			104: begin
				if(in == 0) begin
					state<=105;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=4003;
					out<=10;
				end
				if(in == 3) begin
					state<=2103;
					out<=11;
				end
				if(in == 4) begin
					state<=5992;
					out<=12;
				end
			end
			105: begin
				if(in == 0) begin
					state<=106;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=4004;
					out<=15;
				end
				if(in == 3) begin
					state<=2104;
					out<=16;
				end
				if(in == 4) begin
					state<=5993;
					out<=17;
				end
			end
			106: begin
				if(in == 0) begin
					state<=107;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=4005;
					out<=20;
				end
				if(in == 3) begin
					state<=2105;
					out<=21;
				end
				if(in == 4) begin
					state<=5994;
					out<=22;
				end
			end
			107: begin
				if(in == 0) begin
					state<=108;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=4006;
					out<=25;
				end
				if(in == 3) begin
					state<=2106;
					out<=26;
				end
				if(in == 4) begin
					state<=5995;
					out<=27;
				end
			end
			108: begin
				if(in == 0) begin
					state<=109;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=4007;
					out<=30;
				end
				if(in == 3) begin
					state<=2107;
					out<=31;
				end
				if(in == 4) begin
					state<=5996;
					out<=32;
				end
			end
			109: begin
				if(in == 0) begin
					state<=110;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=4008;
					out<=35;
				end
				if(in == 3) begin
					state<=2108;
					out<=36;
				end
				if(in == 4) begin
					state<=5997;
					out<=37;
				end
			end
			110: begin
				if(in == 0) begin
					state<=111;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=4009;
					out<=40;
				end
				if(in == 3) begin
					state<=2109;
					out<=41;
				end
				if(in == 4) begin
					state<=5998;
					out<=42;
				end
			end
			111: begin
				if(in == 0) begin
					state<=112;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=4010;
					out<=45;
				end
				if(in == 3) begin
					state<=2110;
					out<=46;
				end
				if(in == 4) begin
					state<=5999;
					out<=47;
				end
			end
			112: begin
				if(in == 0) begin
					state<=113;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=4011;
					out<=50;
				end
				if(in == 3) begin
					state<=2111;
					out<=51;
				end
				if(in == 4) begin
					state<=6000;
					out<=52;
				end
			end
			113: begin
				if(in == 0) begin
					state<=114;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=4012;
					out<=55;
				end
				if(in == 3) begin
					state<=2112;
					out<=56;
				end
				if(in == 4) begin
					state<=6001;
					out<=57;
				end
			end
			114: begin
				if(in == 0) begin
					state<=115;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=4013;
					out<=60;
				end
				if(in == 3) begin
					state<=2113;
					out<=61;
				end
				if(in == 4) begin
					state<=6002;
					out<=62;
				end
			end
			115: begin
				if(in == 0) begin
					state<=116;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=4014;
					out<=65;
				end
				if(in == 3) begin
					state<=2114;
					out<=66;
				end
				if(in == 4) begin
					state<=6003;
					out<=67;
				end
			end
			116: begin
				if(in == 0) begin
					state<=117;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=4015;
					out<=70;
				end
				if(in == 3) begin
					state<=2115;
					out<=71;
				end
				if(in == 4) begin
					state<=6004;
					out<=72;
				end
			end
			117: begin
				if(in == 0) begin
					state<=118;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=4016;
					out<=75;
				end
				if(in == 3) begin
					state<=2116;
					out<=76;
				end
				if(in == 4) begin
					state<=6005;
					out<=77;
				end
			end
			118: begin
				if(in == 0) begin
					state<=119;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=4017;
					out<=80;
				end
				if(in == 3) begin
					state<=2117;
					out<=81;
				end
				if(in == 4) begin
					state<=6006;
					out<=82;
				end
			end
			119: begin
				if(in == 0) begin
					state<=1360;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=5249;
					out<=85;
				end
				if(in == 3) begin
					state<=3292;
					out<=86;
				end
				if(in == 4) begin
					state<=7181;
					out<=87;
				end
			end
			120: begin
				if(in == 0) begin
					state<=121;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=4019;
					out<=90;
				end
				if(in == 3) begin
					state<=2119;
					out<=91;
				end
				if(in == 4) begin
					state<=6008;
					out<=92;
				end
			end
			121: begin
				if(in == 0) begin
					state<=122;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=4020;
					out<=95;
				end
				if(in == 3) begin
					state<=2120;
					out<=96;
				end
				if(in == 4) begin
					state<=6009;
					out<=97;
				end
			end
			122: begin
				if(in == 0) begin
					state<=123;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=4021;
					out<=100;
				end
				if(in == 3) begin
					state<=2121;
					out<=101;
				end
				if(in == 4) begin
					state<=6010;
					out<=102;
				end
			end
			123: begin
				if(in == 0) begin
					state<=124;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=4022;
					out<=105;
				end
				if(in == 3) begin
					state<=2122;
					out<=106;
				end
				if(in == 4) begin
					state<=6011;
					out<=107;
				end
			end
			124: begin
				if(in == 0) begin
					state<=125;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=4023;
					out<=110;
				end
				if(in == 3) begin
					state<=2123;
					out<=111;
				end
				if(in == 4) begin
					state<=6012;
					out<=112;
				end
			end
			125: begin
				if(in == 0) begin
					state<=126;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=4024;
					out<=115;
				end
				if(in == 3) begin
					state<=2124;
					out<=116;
				end
				if(in == 4) begin
					state<=6013;
					out<=117;
				end
			end
			126: begin
				if(in == 0) begin
					state<=127;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=4025;
					out<=120;
				end
				if(in == 3) begin
					state<=2125;
					out<=121;
				end
				if(in == 4) begin
					state<=6014;
					out<=122;
				end
			end
			127: begin
				if(in == 0) begin
					state<=128;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=4026;
					out<=125;
				end
				if(in == 3) begin
					state<=2126;
					out<=126;
				end
				if(in == 4) begin
					state<=6015;
					out<=127;
				end
			end
			128: begin
				if(in == 0) begin
					state<=129;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=4027;
					out<=130;
				end
				if(in == 3) begin
					state<=2127;
					out<=131;
				end
				if(in == 4) begin
					state<=6016;
					out<=132;
				end
			end
			129: begin
				if(in == 0) begin
					state<=130;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=4028;
					out<=135;
				end
				if(in == 3) begin
					state<=2128;
					out<=136;
				end
				if(in == 4) begin
					state<=6017;
					out<=137;
				end
			end
			130: begin
				if(in == 0) begin
					state<=131;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=4029;
					out<=140;
				end
				if(in == 3) begin
					state<=2129;
					out<=141;
				end
				if(in == 4) begin
					state<=6018;
					out<=142;
				end
			end
			131: begin
				if(in == 0) begin
					state<=132;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=4030;
					out<=145;
				end
				if(in == 3) begin
					state<=2130;
					out<=146;
				end
				if(in == 4) begin
					state<=6019;
					out<=147;
				end
			end
			132: begin
				if(in == 0) begin
					state<=133;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=4031;
					out<=150;
				end
				if(in == 3) begin
					state<=2131;
					out<=151;
				end
				if(in == 4) begin
					state<=6020;
					out<=152;
				end
			end
			133: begin
				if(in == 0) begin
					state<=134;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=4032;
					out<=155;
				end
				if(in == 3) begin
					state<=2132;
					out<=156;
				end
				if(in == 4) begin
					state<=6021;
					out<=157;
				end
			end
			134: begin
				if(in == 0) begin
					state<=135;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=4033;
					out<=160;
				end
				if(in == 3) begin
					state<=2133;
					out<=161;
				end
				if(in == 4) begin
					state<=6022;
					out<=162;
				end
			end
			135: begin
				if(in == 0) begin
					state<=136;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=4034;
					out<=165;
				end
				if(in == 3) begin
					state<=2134;
					out<=166;
				end
				if(in == 4) begin
					state<=6023;
					out<=167;
				end
			end
			136: begin
				if(in == 0) begin
					state<=137;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=4035;
					out<=170;
				end
				if(in == 3) begin
					state<=2135;
					out<=171;
				end
				if(in == 4) begin
					state<=6024;
					out<=172;
				end
			end
			137: begin
				if(in == 0) begin
					state<=138;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=4036;
					out<=175;
				end
				if(in == 3) begin
					state<=2136;
					out<=176;
				end
				if(in == 4) begin
					state<=6025;
					out<=177;
				end
			end
			138: begin
				if(in == 0) begin
					state<=139;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=4037;
					out<=180;
				end
				if(in == 3) begin
					state<=2137;
					out<=181;
				end
				if(in == 4) begin
					state<=6026;
					out<=182;
				end
			end
			139: begin
				if(in == 0) begin
					state<=140;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=4038;
					out<=185;
				end
				if(in == 3) begin
					state<=2138;
					out<=186;
				end
				if(in == 4) begin
					state<=6027;
					out<=187;
				end
			end
			140: begin
				if(in == 0) begin
					state<=141;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=4039;
					out<=190;
				end
				if(in == 3) begin
					state<=2139;
					out<=191;
				end
				if(in == 4) begin
					state<=6028;
					out<=192;
				end
			end
			141: begin
				if(in == 0) begin
					state<=142;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=4040;
					out<=195;
				end
				if(in == 3) begin
					state<=2140;
					out<=196;
				end
				if(in == 4) begin
					state<=6029;
					out<=197;
				end
			end
			142: begin
				if(in == 0) begin
					state<=143;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=4041;
					out<=200;
				end
				if(in == 3) begin
					state<=2141;
					out<=201;
				end
				if(in == 4) begin
					state<=6030;
					out<=202;
				end
			end
			143: begin
				if(in == 0) begin
					state<=144;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=4042;
					out<=205;
				end
				if(in == 3) begin
					state<=2142;
					out<=206;
				end
				if(in == 4) begin
					state<=6031;
					out<=207;
				end
			end
			144: begin
				if(in == 0) begin
					state<=145;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=4043;
					out<=210;
				end
				if(in == 3) begin
					state<=2143;
					out<=211;
				end
				if(in == 4) begin
					state<=6032;
					out<=212;
				end
			end
			145: begin
				if(in == 0) begin
					state<=146;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=4044;
					out<=215;
				end
				if(in == 3) begin
					state<=2144;
					out<=216;
				end
				if(in == 4) begin
					state<=6033;
					out<=217;
				end
			end
			146: begin
				if(in == 0) begin
					state<=147;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=4045;
					out<=220;
				end
				if(in == 3) begin
					state<=2145;
					out<=221;
				end
				if(in == 4) begin
					state<=6034;
					out<=222;
				end
			end
			147: begin
				if(in == 0) begin
					state<=148;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=4046;
					out<=225;
				end
				if(in == 3) begin
					state<=2146;
					out<=226;
				end
				if(in == 4) begin
					state<=6035;
					out<=227;
				end
			end
			148: begin
				if(in == 0) begin
					state<=149;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=4047;
					out<=230;
				end
				if(in == 3) begin
					state<=2147;
					out<=231;
				end
				if(in == 4) begin
					state<=6036;
					out<=232;
				end
			end
			149: begin
				if(in == 0) begin
					state<=150;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=4048;
					out<=235;
				end
				if(in == 3) begin
					state<=2148;
					out<=236;
				end
				if(in == 4) begin
					state<=6037;
					out<=237;
				end
			end
			150: begin
				if(in == 0) begin
					state<=151;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=4049;
					out<=240;
				end
				if(in == 3) begin
					state<=2149;
					out<=241;
				end
				if(in == 4) begin
					state<=6038;
					out<=242;
				end
			end
			151: begin
				if(in == 0) begin
					state<=152;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=4050;
					out<=245;
				end
				if(in == 3) begin
					state<=2150;
					out<=246;
				end
				if(in == 4) begin
					state<=6039;
					out<=247;
				end
			end
			152: begin
				if(in == 0) begin
					state<=153;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=4051;
					out<=250;
				end
				if(in == 3) begin
					state<=2151;
					out<=251;
				end
				if(in == 4) begin
					state<=6040;
					out<=252;
				end
			end
			153: begin
				if(in == 0) begin
					state<=154;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=4052;
					out<=255;
				end
				if(in == 3) begin
					state<=2152;
					out<=0;
				end
				if(in == 4) begin
					state<=6041;
					out<=1;
				end
			end
			154: begin
				if(in == 0) begin
					state<=155;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=4053;
					out<=4;
				end
				if(in == 3) begin
					state<=2153;
					out<=5;
				end
				if(in == 4) begin
					state<=6042;
					out<=6;
				end
			end
			155: begin
				if(in == 0) begin
					state<=156;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=4054;
					out<=9;
				end
				if(in == 3) begin
					state<=2154;
					out<=10;
				end
				if(in == 4) begin
					state<=6043;
					out<=11;
				end
			end
			156: begin
				if(in == 0) begin
					state<=157;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=4055;
					out<=14;
				end
				if(in == 3) begin
					state<=2155;
					out<=15;
				end
				if(in == 4) begin
					state<=6044;
					out<=16;
				end
			end
			157: begin
				if(in == 0) begin
					state<=158;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=4056;
					out<=19;
				end
				if(in == 3) begin
					state<=2156;
					out<=20;
				end
				if(in == 4) begin
					state<=6045;
					out<=21;
				end
			end
			158: begin
				if(in == 0) begin
					state<=159;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=4057;
					out<=24;
				end
				if(in == 3) begin
					state<=2157;
					out<=25;
				end
				if(in == 4) begin
					state<=6046;
					out<=26;
				end
			end
			159: begin
				if(in == 0) begin
					state<=160;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=4058;
					out<=29;
				end
				if(in == 3) begin
					state<=2158;
					out<=30;
				end
				if(in == 4) begin
					state<=6047;
					out<=31;
				end
			end
			160: begin
				if(in == 0) begin
					state<=161;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=4059;
					out<=34;
				end
				if(in == 3) begin
					state<=2159;
					out<=35;
				end
				if(in == 4) begin
					state<=6048;
					out<=36;
				end
			end
			161: begin
				if(in == 0) begin
					state<=162;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=4060;
					out<=39;
				end
				if(in == 3) begin
					state<=2160;
					out<=40;
				end
				if(in == 4) begin
					state<=6049;
					out<=41;
				end
			end
			162: begin
				if(in == 0) begin
					state<=163;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=4061;
					out<=44;
				end
				if(in == 3) begin
					state<=2161;
					out<=45;
				end
				if(in == 4) begin
					state<=6050;
					out<=46;
				end
			end
			163: begin
				if(in == 0) begin
					state<=164;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=4062;
					out<=49;
				end
				if(in == 3) begin
					state<=2162;
					out<=50;
				end
				if(in == 4) begin
					state<=6051;
					out<=51;
				end
			end
			164: begin
				if(in == 0) begin
					state<=165;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=4063;
					out<=54;
				end
				if(in == 3) begin
					state<=2163;
					out<=55;
				end
				if(in == 4) begin
					state<=6052;
					out<=56;
				end
			end
			165: begin
				if(in == 0) begin
					state<=166;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=4064;
					out<=59;
				end
				if(in == 3) begin
					state<=2164;
					out<=60;
				end
				if(in == 4) begin
					state<=6053;
					out<=61;
				end
			end
			166: begin
				if(in == 0) begin
					state<=167;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=4065;
					out<=64;
				end
				if(in == 3) begin
					state<=2165;
					out<=65;
				end
				if(in == 4) begin
					state<=6054;
					out<=66;
				end
			end
			167: begin
				if(in == 0) begin
					state<=168;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=4066;
					out<=69;
				end
				if(in == 3) begin
					state<=2166;
					out<=70;
				end
				if(in == 4) begin
					state<=6055;
					out<=71;
				end
			end
			168: begin
				if(in == 0) begin
					state<=169;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=4067;
					out<=74;
				end
				if(in == 3) begin
					state<=2167;
					out<=75;
				end
				if(in == 4) begin
					state<=6056;
					out<=76;
				end
			end
			169: begin
				if(in == 0) begin
					state<=170;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=4068;
					out<=79;
				end
				if(in == 3) begin
					state<=2168;
					out<=80;
				end
				if(in == 4) begin
					state<=6057;
					out<=81;
				end
			end
			170: begin
				if(in == 0) begin
					state<=171;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=4069;
					out<=84;
				end
				if(in == 3) begin
					state<=2169;
					out<=85;
				end
				if(in == 4) begin
					state<=6058;
					out<=86;
				end
			end
			171: begin
				if(in == 0) begin
					state<=172;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=4070;
					out<=89;
				end
				if(in == 3) begin
					state<=2170;
					out<=90;
				end
				if(in == 4) begin
					state<=6059;
					out<=91;
				end
			end
			172: begin
				if(in == 0) begin
					state<=173;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=4071;
					out<=94;
				end
				if(in == 3) begin
					state<=2171;
					out<=95;
				end
				if(in == 4) begin
					state<=6060;
					out<=96;
				end
			end
			173: begin
				if(in == 0) begin
					state<=174;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=4072;
					out<=99;
				end
				if(in == 3) begin
					state<=2172;
					out<=100;
				end
				if(in == 4) begin
					state<=6061;
					out<=101;
				end
			end
			174: begin
				if(in == 0) begin
					state<=175;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=4073;
					out<=104;
				end
				if(in == 3) begin
					state<=2173;
					out<=105;
				end
				if(in == 4) begin
					state<=6062;
					out<=106;
				end
			end
			175: begin
				if(in == 0) begin
					state<=176;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=4074;
					out<=109;
				end
				if(in == 3) begin
					state<=2174;
					out<=110;
				end
				if(in == 4) begin
					state<=6063;
					out<=111;
				end
			end
			176: begin
				if(in == 0) begin
					state<=177;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=4075;
					out<=114;
				end
				if(in == 3) begin
					state<=2175;
					out<=115;
				end
				if(in == 4) begin
					state<=6064;
					out<=116;
				end
			end
			177: begin
				if(in == 0) begin
					state<=178;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=4076;
					out<=119;
				end
				if(in == 3) begin
					state<=2176;
					out<=120;
				end
				if(in == 4) begin
					state<=6065;
					out<=121;
				end
			end
			178: begin
				if(in == 0) begin
					state<=179;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=4077;
					out<=124;
				end
				if(in == 3) begin
					state<=2177;
					out<=125;
				end
				if(in == 4) begin
					state<=6066;
					out<=126;
				end
			end
			179: begin
				if(in == 0) begin
					state<=180;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=4078;
					out<=129;
				end
				if(in == 3) begin
					state<=2178;
					out<=130;
				end
				if(in == 4) begin
					state<=6067;
					out<=131;
				end
			end
			180: begin
				if(in == 0) begin
					state<=181;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=4079;
					out<=134;
				end
				if(in == 3) begin
					state<=2179;
					out<=135;
				end
				if(in == 4) begin
					state<=6068;
					out<=136;
				end
			end
			181: begin
				if(in == 0) begin
					state<=182;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=4080;
					out<=139;
				end
				if(in == 3) begin
					state<=2180;
					out<=140;
				end
				if(in == 4) begin
					state<=6069;
					out<=141;
				end
			end
			182: begin
				if(in == 0) begin
					state<=183;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=4081;
					out<=144;
				end
				if(in == 3) begin
					state<=2181;
					out<=145;
				end
				if(in == 4) begin
					state<=6070;
					out<=146;
				end
			end
			183: begin
				if(in == 0) begin
					state<=184;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=4082;
					out<=149;
				end
				if(in == 3) begin
					state<=2182;
					out<=150;
				end
				if(in == 4) begin
					state<=6071;
					out<=151;
				end
			end
			184: begin
				if(in == 0) begin
					state<=185;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=4083;
					out<=154;
				end
				if(in == 3) begin
					state<=2183;
					out<=155;
				end
				if(in == 4) begin
					state<=6072;
					out<=156;
				end
			end
			185: begin
				if(in == 0) begin
					state<=186;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=4084;
					out<=159;
				end
				if(in == 3) begin
					state<=2184;
					out<=160;
				end
				if(in == 4) begin
					state<=6073;
					out<=161;
				end
			end
			186: begin
				if(in == 0) begin
					state<=187;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=4085;
					out<=164;
				end
				if(in == 3) begin
					state<=2185;
					out<=165;
				end
				if(in == 4) begin
					state<=6074;
					out<=166;
				end
			end
			187: begin
				if(in == 0) begin
					state<=188;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=4086;
					out<=169;
				end
				if(in == 3) begin
					state<=2186;
					out<=170;
				end
				if(in == 4) begin
					state<=6075;
					out<=171;
				end
			end
			188: begin
				if(in == 0) begin
					state<=1391;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=5280;
					out<=174;
				end
				if(in == 3) begin
					state<=3323;
					out<=175;
				end
				if(in == 4) begin
					state<=7212;
					out<=176;
				end
			end
			189: begin
				if(in == 0) begin
					state<=190;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=4088;
					out<=179;
				end
				if(in == 3) begin
					state<=2188;
					out<=180;
				end
				if(in == 4) begin
					state<=6077;
					out<=181;
				end
			end
			190: begin
				if(in == 0) begin
					state<=191;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=4089;
					out<=184;
				end
				if(in == 3) begin
					state<=2189;
					out<=185;
				end
				if(in == 4) begin
					state<=6078;
					out<=186;
				end
			end
			191: begin
				if(in == 0) begin
					state<=192;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=4090;
					out<=189;
				end
				if(in == 3) begin
					state<=2190;
					out<=190;
				end
				if(in == 4) begin
					state<=6079;
					out<=191;
				end
			end
			192: begin
				if(in == 0) begin
					state<=193;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=4091;
					out<=194;
				end
				if(in == 3) begin
					state<=2191;
					out<=195;
				end
				if(in == 4) begin
					state<=6080;
					out<=196;
				end
			end
			193: begin
				if(in == 0) begin
					state<=194;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=4092;
					out<=199;
				end
				if(in == 3) begin
					state<=2192;
					out<=200;
				end
				if(in == 4) begin
					state<=6081;
					out<=201;
				end
			end
			194: begin
				if(in == 0) begin
					state<=195;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=4093;
					out<=204;
				end
				if(in == 3) begin
					state<=2193;
					out<=205;
				end
				if(in == 4) begin
					state<=6082;
					out<=206;
				end
			end
			195: begin
				if(in == 0) begin
					state<=196;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=4094;
					out<=209;
				end
				if(in == 3) begin
					state<=2194;
					out<=210;
				end
				if(in == 4) begin
					state<=6083;
					out<=211;
				end
			end
			196: begin
				if(in == 0) begin
					state<=197;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=4095;
					out<=214;
				end
				if(in == 3) begin
					state<=2195;
					out<=215;
				end
				if(in == 4) begin
					state<=6084;
					out<=216;
				end
			end
			197: begin
				if(in == 0) begin
					state<=198;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=4096;
					out<=219;
				end
				if(in == 3) begin
					state<=2196;
					out<=220;
				end
				if(in == 4) begin
					state<=6085;
					out<=221;
				end
			end
			198: begin
				if(in == 0) begin
					state<=199;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=4097;
					out<=224;
				end
				if(in == 3) begin
					state<=2197;
					out<=225;
				end
				if(in == 4) begin
					state<=6086;
					out<=226;
				end
			end
			199: begin
				if(in == 0) begin
					state<=200;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=4098;
					out<=229;
				end
				if(in == 3) begin
					state<=2198;
					out<=230;
				end
				if(in == 4) begin
					state<=6087;
					out<=231;
				end
			end
			200: begin
				if(in == 0) begin
					state<=201;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=4099;
					out<=234;
				end
				if(in == 3) begin
					state<=2199;
					out<=235;
				end
				if(in == 4) begin
					state<=6088;
					out<=236;
				end
			end
			201: begin
				if(in == 0) begin
					state<=202;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=4100;
					out<=239;
				end
				if(in == 3) begin
					state<=2200;
					out<=240;
				end
				if(in == 4) begin
					state<=6089;
					out<=241;
				end
			end
			202: begin
				if(in == 0) begin
					state<=203;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=4101;
					out<=244;
				end
				if(in == 3) begin
					state<=2201;
					out<=245;
				end
				if(in == 4) begin
					state<=6090;
					out<=246;
				end
			end
			203: begin
				if(in == 0) begin
					state<=204;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=4102;
					out<=249;
				end
				if(in == 3) begin
					state<=2202;
					out<=250;
				end
				if(in == 4) begin
					state<=6091;
					out<=251;
				end
			end
			204: begin
				if(in == 0) begin
					state<=205;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=4103;
					out<=254;
				end
				if(in == 3) begin
					state<=2203;
					out<=255;
				end
				if(in == 4) begin
					state<=6092;
					out<=0;
				end
			end
			205: begin
				if(in == 0) begin
					state<=206;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=4104;
					out<=3;
				end
				if(in == 3) begin
					state<=2204;
					out<=4;
				end
				if(in == 4) begin
					state<=6093;
					out<=5;
				end
			end
			206: begin
				if(in == 0) begin
					state<=207;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=4105;
					out<=8;
				end
				if(in == 3) begin
					state<=2205;
					out<=9;
				end
				if(in == 4) begin
					state<=6094;
					out<=10;
				end
			end
			207: begin
				if(in == 0) begin
					state<=208;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=4106;
					out<=13;
				end
				if(in == 3) begin
					state<=2206;
					out<=14;
				end
				if(in == 4) begin
					state<=6095;
					out<=15;
				end
			end
			208: begin
				if(in == 0) begin
					state<=209;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=4107;
					out<=18;
				end
				if(in == 3) begin
					state<=2207;
					out<=19;
				end
				if(in == 4) begin
					state<=6096;
					out<=20;
				end
			end
			209: begin
				if(in == 0) begin
					state<=210;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=4108;
					out<=23;
				end
				if(in == 3) begin
					state<=2208;
					out<=24;
				end
				if(in == 4) begin
					state<=6097;
					out<=25;
				end
			end
			210: begin
				if(in == 0) begin
					state<=211;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=4109;
					out<=28;
				end
				if(in == 3) begin
					state<=2209;
					out<=29;
				end
				if(in == 4) begin
					state<=6098;
					out<=30;
				end
			end
			211: begin
				if(in == 0) begin
					state<=212;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=4110;
					out<=33;
				end
				if(in == 3) begin
					state<=2210;
					out<=34;
				end
				if(in == 4) begin
					state<=6099;
					out<=35;
				end
			end
			212: begin
				if(in == 0) begin
					state<=213;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=4111;
					out<=38;
				end
				if(in == 3) begin
					state<=2211;
					out<=39;
				end
				if(in == 4) begin
					state<=6100;
					out<=40;
				end
			end
			213: begin
				if(in == 0) begin
					state<=214;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=4112;
					out<=43;
				end
				if(in == 3) begin
					state<=2212;
					out<=44;
				end
				if(in == 4) begin
					state<=6101;
					out<=45;
				end
			end
			214: begin
				if(in == 0) begin
					state<=215;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=4113;
					out<=48;
				end
				if(in == 3) begin
					state<=2213;
					out<=49;
				end
				if(in == 4) begin
					state<=6102;
					out<=50;
				end
			end
			215: begin
				if(in == 0) begin
					state<=216;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=4114;
					out<=53;
				end
				if(in == 3) begin
					state<=2214;
					out<=54;
				end
				if(in == 4) begin
					state<=6103;
					out<=55;
				end
			end
			216: begin
				if(in == 0) begin
					state<=217;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=4115;
					out<=58;
				end
				if(in == 3) begin
					state<=2215;
					out<=59;
				end
				if(in == 4) begin
					state<=6104;
					out<=60;
				end
			end
			217: begin
				if(in == 0) begin
					state<=218;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=4116;
					out<=63;
				end
				if(in == 3) begin
					state<=2216;
					out<=64;
				end
				if(in == 4) begin
					state<=6105;
					out<=65;
				end
			end
			218: begin
				if(in == 0) begin
					state<=219;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=4117;
					out<=68;
				end
				if(in == 3) begin
					state<=2217;
					out<=69;
				end
				if(in == 4) begin
					state<=6106;
					out<=70;
				end
			end
			219: begin
				if(in == 0) begin
					state<=220;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=4118;
					out<=73;
				end
				if(in == 3) begin
					state<=2218;
					out<=74;
				end
				if(in == 4) begin
					state<=6107;
					out<=75;
				end
			end
			220: begin
				if(in == 0) begin
					state<=221;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=4119;
					out<=78;
				end
				if(in == 3) begin
					state<=2219;
					out<=79;
				end
				if(in == 4) begin
					state<=6108;
					out<=80;
				end
			end
			221: begin
				if(in == 0) begin
					state<=222;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=4120;
					out<=83;
				end
				if(in == 3) begin
					state<=2220;
					out<=84;
				end
				if(in == 4) begin
					state<=6109;
					out<=85;
				end
			end
			222: begin
				if(in == 0) begin
					state<=223;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=4121;
					out<=88;
				end
				if(in == 3) begin
					state<=2221;
					out<=89;
				end
				if(in == 4) begin
					state<=6110;
					out<=90;
				end
			end
			223: begin
				if(in == 0) begin
					state<=224;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=4122;
					out<=93;
				end
				if(in == 3) begin
					state<=2222;
					out<=94;
				end
				if(in == 4) begin
					state<=6111;
					out<=95;
				end
			end
			224: begin
				if(in == 0) begin
					state<=225;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=4123;
					out<=98;
				end
				if(in == 3) begin
					state<=2223;
					out<=99;
				end
				if(in == 4) begin
					state<=6112;
					out<=100;
				end
			end
			225: begin
				if(in == 0) begin
					state<=226;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=4124;
					out<=103;
				end
				if(in == 3) begin
					state<=2224;
					out<=104;
				end
				if(in == 4) begin
					state<=6113;
					out<=105;
				end
			end
			226: begin
				if(in == 0) begin
					state<=227;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=4125;
					out<=108;
				end
				if(in == 3) begin
					state<=2225;
					out<=109;
				end
				if(in == 4) begin
					state<=6114;
					out<=110;
				end
			end
			227: begin
				if(in == 0) begin
					state<=228;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=4126;
					out<=113;
				end
				if(in == 3) begin
					state<=2226;
					out<=114;
				end
				if(in == 4) begin
					state<=6115;
					out<=115;
				end
			end
			228: begin
				if(in == 0) begin
					state<=229;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=4127;
					out<=118;
				end
				if(in == 3) begin
					state<=2227;
					out<=119;
				end
				if(in == 4) begin
					state<=6116;
					out<=120;
				end
			end
			229: begin
				if(in == 0) begin
					state<=230;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=4128;
					out<=123;
				end
				if(in == 3) begin
					state<=2228;
					out<=124;
				end
				if(in == 4) begin
					state<=6117;
					out<=125;
				end
			end
			230: begin
				if(in == 0) begin
					state<=231;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=4129;
					out<=128;
				end
				if(in == 3) begin
					state<=2229;
					out<=129;
				end
				if(in == 4) begin
					state<=6118;
					out<=130;
				end
			end
			231: begin
				if(in == 0) begin
					state<=232;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=4130;
					out<=133;
				end
				if(in == 3) begin
					state<=2230;
					out<=134;
				end
				if(in == 4) begin
					state<=6119;
					out<=135;
				end
			end
			232: begin
				if(in == 0) begin
					state<=233;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=4131;
					out<=138;
				end
				if(in == 3) begin
					state<=2231;
					out<=139;
				end
				if(in == 4) begin
					state<=6120;
					out<=140;
				end
			end
			233: begin
				if(in == 0) begin
					state<=234;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=4132;
					out<=143;
				end
				if(in == 3) begin
					state<=2232;
					out<=144;
				end
				if(in == 4) begin
					state<=6121;
					out<=145;
				end
			end
			234: begin
				if(in == 0) begin
					state<=235;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=4133;
					out<=148;
				end
				if(in == 3) begin
					state<=2233;
					out<=149;
				end
				if(in == 4) begin
					state<=6122;
					out<=150;
				end
			end
			235: begin
				if(in == 0) begin
					state<=236;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=4134;
					out<=153;
				end
				if(in == 3) begin
					state<=2234;
					out<=154;
				end
				if(in == 4) begin
					state<=6123;
					out<=155;
				end
			end
			236: begin
				if(in == 0) begin
					state<=237;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=4135;
					out<=158;
				end
				if(in == 3) begin
					state<=2235;
					out<=159;
				end
				if(in == 4) begin
					state<=6124;
					out<=160;
				end
			end
			237: begin
				if(in == 0) begin
					state<=238;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=4136;
					out<=163;
				end
				if(in == 3) begin
					state<=2236;
					out<=164;
				end
				if(in == 4) begin
					state<=6125;
					out<=165;
				end
			end
			238: begin
				if(in == 0) begin
					state<=239;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=4137;
					out<=168;
				end
				if(in == 3) begin
					state<=2237;
					out<=169;
				end
				if(in == 4) begin
					state<=6126;
					out<=170;
				end
			end
			239: begin
				if(in == 0) begin
					state<=240;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=4138;
					out<=173;
				end
				if(in == 3) begin
					state<=2238;
					out<=174;
				end
				if(in == 4) begin
					state<=6127;
					out<=175;
				end
			end
			240: begin
				if(in == 0) begin
					state<=241;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=4139;
					out<=178;
				end
				if(in == 3) begin
					state<=2239;
					out<=179;
				end
				if(in == 4) begin
					state<=6128;
					out<=180;
				end
			end
			241: begin
				if(in == 0) begin
					state<=242;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=4140;
					out<=183;
				end
				if(in == 3) begin
					state<=2240;
					out<=184;
				end
				if(in == 4) begin
					state<=6129;
					out<=185;
				end
			end
			242: begin
				if(in == 0) begin
					state<=243;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=4141;
					out<=188;
				end
				if(in == 3) begin
					state<=2241;
					out<=189;
				end
				if(in == 4) begin
					state<=6130;
					out<=190;
				end
			end
			243: begin
				if(in == 0) begin
					state<=244;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=4142;
					out<=193;
				end
				if(in == 3) begin
					state<=2242;
					out<=194;
				end
				if(in == 4) begin
					state<=6131;
					out<=195;
				end
			end
			244: begin
				if(in == 0) begin
					state<=245;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=4143;
					out<=198;
				end
				if(in == 3) begin
					state<=2243;
					out<=199;
				end
				if(in == 4) begin
					state<=6132;
					out<=200;
				end
			end
			245: begin
				if(in == 0) begin
					state<=246;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=4144;
					out<=203;
				end
				if(in == 3) begin
					state<=2244;
					out<=204;
				end
				if(in == 4) begin
					state<=6133;
					out<=205;
				end
			end
			246: begin
				if(in == 0) begin
					state<=247;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=4145;
					out<=208;
				end
				if(in == 3) begin
					state<=2245;
					out<=209;
				end
				if(in == 4) begin
					state<=6134;
					out<=210;
				end
			end
			247: begin
				if(in == 0) begin
					state<=248;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=4146;
					out<=213;
				end
				if(in == 3) begin
					state<=2246;
					out<=214;
				end
				if(in == 4) begin
					state<=6135;
					out<=215;
				end
			end
			248: begin
				if(in == 0) begin
					state<=249;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=4147;
					out<=218;
				end
				if(in == 3) begin
					state<=2247;
					out<=219;
				end
				if(in == 4) begin
					state<=6136;
					out<=220;
				end
			end
			249: begin
				if(in == 0) begin
					state<=250;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=4148;
					out<=223;
				end
				if(in == 3) begin
					state<=2248;
					out<=224;
				end
				if(in == 4) begin
					state<=6137;
					out<=225;
				end
			end
			250: begin
				if(in == 0) begin
					state<=251;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=4149;
					out<=228;
				end
				if(in == 3) begin
					state<=2249;
					out<=229;
				end
				if(in == 4) begin
					state<=6138;
					out<=230;
				end
			end
			251: begin
				if(in == 0) begin
					state<=252;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=4150;
					out<=233;
				end
				if(in == 3) begin
					state<=2250;
					out<=234;
				end
				if(in == 4) begin
					state<=6139;
					out<=235;
				end
			end
			252: begin
				if(in == 0) begin
					state<=253;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=4151;
					out<=238;
				end
				if(in == 3) begin
					state<=2251;
					out<=239;
				end
				if(in == 4) begin
					state<=6140;
					out<=240;
				end
			end
			253: begin
				if(in == 0) begin
					state<=254;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=4152;
					out<=243;
				end
				if(in == 3) begin
					state<=2252;
					out<=244;
				end
				if(in == 4) begin
					state<=6141;
					out<=245;
				end
			end
			254: begin
				if(in == 0) begin
					state<=255;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=4153;
					out<=248;
				end
				if(in == 3) begin
					state<=2253;
					out<=249;
				end
				if(in == 4) begin
					state<=6142;
					out<=250;
				end
			end
			255: begin
				if(in == 0) begin
					state<=256;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=4154;
					out<=253;
				end
				if(in == 3) begin
					state<=2254;
					out<=254;
				end
				if(in == 4) begin
					state<=6143;
					out<=255;
				end
			end
			256: begin
				if(in == 0) begin
					state<=257;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=4155;
					out<=2;
				end
				if(in == 3) begin
					state<=2255;
					out<=3;
				end
				if(in == 4) begin
					state<=6144;
					out<=4;
				end
			end
			257: begin
				if(in == 0) begin
					state<=1422;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=5311;
					out<=7;
				end
				if(in == 3) begin
					state<=3354;
					out<=8;
				end
				if(in == 4) begin
					state<=7243;
					out<=9;
				end
			end
			258: begin
				if(in == 0) begin
					state<=259;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=4157;
					out<=12;
				end
				if(in == 3) begin
					state<=2257;
					out<=13;
				end
				if(in == 4) begin
					state<=6146;
					out<=14;
				end
			end
			259: begin
				if(in == 0) begin
					state<=260;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=4158;
					out<=17;
				end
				if(in == 3) begin
					state<=2258;
					out<=18;
				end
				if(in == 4) begin
					state<=6147;
					out<=19;
				end
			end
			260: begin
				if(in == 0) begin
					state<=261;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=4159;
					out<=22;
				end
				if(in == 3) begin
					state<=2259;
					out<=23;
				end
				if(in == 4) begin
					state<=6148;
					out<=24;
				end
			end
			261: begin
				if(in == 0) begin
					state<=262;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=4160;
					out<=27;
				end
				if(in == 3) begin
					state<=2260;
					out<=28;
				end
				if(in == 4) begin
					state<=6149;
					out<=29;
				end
			end
			262: begin
				if(in == 0) begin
					state<=263;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=4161;
					out<=32;
				end
				if(in == 3) begin
					state<=2261;
					out<=33;
				end
				if(in == 4) begin
					state<=6150;
					out<=34;
				end
			end
			263: begin
				if(in == 0) begin
					state<=264;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=4162;
					out<=37;
				end
				if(in == 3) begin
					state<=2262;
					out<=38;
				end
				if(in == 4) begin
					state<=6151;
					out<=39;
				end
			end
			264: begin
				if(in == 0) begin
					state<=265;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=4163;
					out<=42;
				end
				if(in == 3) begin
					state<=2263;
					out<=43;
				end
				if(in == 4) begin
					state<=6152;
					out<=44;
				end
			end
			265: begin
				if(in == 0) begin
					state<=266;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=4164;
					out<=47;
				end
				if(in == 3) begin
					state<=2264;
					out<=48;
				end
				if(in == 4) begin
					state<=6153;
					out<=49;
				end
			end
			266: begin
				if(in == 0) begin
					state<=267;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=4165;
					out<=52;
				end
				if(in == 3) begin
					state<=2265;
					out<=53;
				end
				if(in == 4) begin
					state<=6154;
					out<=54;
				end
			end
			267: begin
				if(in == 0) begin
					state<=268;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=4166;
					out<=57;
				end
				if(in == 3) begin
					state<=2266;
					out<=58;
				end
				if(in == 4) begin
					state<=6155;
					out<=59;
				end
			end
			268: begin
				if(in == 0) begin
					state<=269;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=4167;
					out<=62;
				end
				if(in == 3) begin
					state<=2267;
					out<=63;
				end
				if(in == 4) begin
					state<=6156;
					out<=64;
				end
			end
			269: begin
				if(in == 0) begin
					state<=270;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=4168;
					out<=67;
				end
				if(in == 3) begin
					state<=2268;
					out<=68;
				end
				if(in == 4) begin
					state<=6157;
					out<=69;
				end
			end
			270: begin
				if(in == 0) begin
					state<=271;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=4169;
					out<=72;
				end
				if(in == 3) begin
					state<=2269;
					out<=73;
				end
				if(in == 4) begin
					state<=6158;
					out<=74;
				end
			end
			271: begin
				if(in == 0) begin
					state<=272;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=4170;
					out<=77;
				end
				if(in == 3) begin
					state<=2270;
					out<=78;
				end
				if(in == 4) begin
					state<=6159;
					out<=79;
				end
			end
			272: begin
				if(in == 0) begin
					state<=273;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=4171;
					out<=82;
				end
				if(in == 3) begin
					state<=2271;
					out<=83;
				end
				if(in == 4) begin
					state<=6160;
					out<=84;
				end
			end
			273: begin
				if(in == 0) begin
					state<=274;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=4172;
					out<=87;
				end
				if(in == 3) begin
					state<=2272;
					out<=88;
				end
				if(in == 4) begin
					state<=6161;
					out<=89;
				end
			end
			274: begin
				if(in == 0) begin
					state<=275;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=4173;
					out<=92;
				end
				if(in == 3) begin
					state<=2273;
					out<=93;
				end
				if(in == 4) begin
					state<=6162;
					out<=94;
				end
			end
			275: begin
				if(in == 0) begin
					state<=276;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=4174;
					out<=97;
				end
				if(in == 3) begin
					state<=2274;
					out<=98;
				end
				if(in == 4) begin
					state<=6163;
					out<=99;
				end
			end
			276: begin
				if(in == 0) begin
					state<=277;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=4175;
					out<=102;
				end
				if(in == 3) begin
					state<=2275;
					out<=103;
				end
				if(in == 4) begin
					state<=6164;
					out<=104;
				end
			end
			277: begin
				if(in == 0) begin
					state<=278;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=4176;
					out<=107;
				end
				if(in == 3) begin
					state<=2276;
					out<=108;
				end
				if(in == 4) begin
					state<=6165;
					out<=109;
				end
			end
			278: begin
				if(in == 0) begin
					state<=279;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=4177;
					out<=112;
				end
				if(in == 3) begin
					state<=2277;
					out<=113;
				end
				if(in == 4) begin
					state<=6166;
					out<=114;
				end
			end
			279: begin
				if(in == 0) begin
					state<=280;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=4178;
					out<=117;
				end
				if(in == 3) begin
					state<=2278;
					out<=118;
				end
				if(in == 4) begin
					state<=6167;
					out<=119;
				end
			end
			280: begin
				if(in == 0) begin
					state<=281;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=4179;
					out<=122;
				end
				if(in == 3) begin
					state<=2279;
					out<=123;
				end
				if(in == 4) begin
					state<=6168;
					out<=124;
				end
			end
			281: begin
				if(in == 0) begin
					state<=282;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=4180;
					out<=127;
				end
				if(in == 3) begin
					state<=2280;
					out<=128;
				end
				if(in == 4) begin
					state<=6169;
					out<=129;
				end
			end
			282: begin
				if(in == 0) begin
					state<=283;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=4181;
					out<=132;
				end
				if(in == 3) begin
					state<=2281;
					out<=133;
				end
				if(in == 4) begin
					state<=6170;
					out<=134;
				end
			end
			283: begin
				if(in == 0) begin
					state<=284;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=4182;
					out<=137;
				end
				if(in == 3) begin
					state<=2282;
					out<=138;
				end
				if(in == 4) begin
					state<=6171;
					out<=139;
				end
			end
			284: begin
				if(in == 0) begin
					state<=285;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=4183;
					out<=142;
				end
				if(in == 3) begin
					state<=2283;
					out<=143;
				end
				if(in == 4) begin
					state<=6172;
					out<=144;
				end
			end
			285: begin
				if(in == 0) begin
					state<=286;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=4184;
					out<=147;
				end
				if(in == 3) begin
					state<=2284;
					out<=148;
				end
				if(in == 4) begin
					state<=6173;
					out<=149;
				end
			end
			286: begin
				if(in == 0) begin
					state<=287;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=4185;
					out<=152;
				end
				if(in == 3) begin
					state<=2285;
					out<=153;
				end
				if(in == 4) begin
					state<=6174;
					out<=154;
				end
			end
			287: begin
				if(in == 0) begin
					state<=288;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=4186;
					out<=157;
				end
				if(in == 3) begin
					state<=2286;
					out<=158;
				end
				if(in == 4) begin
					state<=6175;
					out<=159;
				end
			end
			288: begin
				if(in == 0) begin
					state<=289;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=4187;
					out<=162;
				end
				if(in == 3) begin
					state<=2287;
					out<=163;
				end
				if(in == 4) begin
					state<=6176;
					out<=164;
				end
			end
			289: begin
				if(in == 0) begin
					state<=290;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=4188;
					out<=167;
				end
				if(in == 3) begin
					state<=2288;
					out<=168;
				end
				if(in == 4) begin
					state<=6177;
					out<=169;
				end
			end
			290: begin
				if(in == 0) begin
					state<=291;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=4189;
					out<=172;
				end
				if(in == 3) begin
					state<=2289;
					out<=173;
				end
				if(in == 4) begin
					state<=6178;
					out<=174;
				end
			end
			291: begin
				if(in == 0) begin
					state<=292;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=4190;
					out<=177;
				end
				if(in == 3) begin
					state<=2290;
					out<=178;
				end
				if(in == 4) begin
					state<=6179;
					out<=179;
				end
			end
			292: begin
				if(in == 0) begin
					state<=293;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=4191;
					out<=182;
				end
				if(in == 3) begin
					state<=2291;
					out<=183;
				end
				if(in == 4) begin
					state<=6180;
					out<=184;
				end
			end
			293: begin
				if(in == 0) begin
					state<=294;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=4192;
					out<=187;
				end
				if(in == 3) begin
					state<=2292;
					out<=188;
				end
				if(in == 4) begin
					state<=6181;
					out<=189;
				end
			end
			294: begin
				if(in == 0) begin
					state<=295;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=4193;
					out<=192;
				end
				if(in == 3) begin
					state<=2293;
					out<=193;
				end
				if(in == 4) begin
					state<=6182;
					out<=194;
				end
			end
			295: begin
				if(in == 0) begin
					state<=296;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=4194;
					out<=197;
				end
				if(in == 3) begin
					state<=2294;
					out<=198;
				end
				if(in == 4) begin
					state<=6183;
					out<=199;
				end
			end
			296: begin
				if(in == 0) begin
					state<=297;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=4195;
					out<=202;
				end
				if(in == 3) begin
					state<=2295;
					out<=203;
				end
				if(in == 4) begin
					state<=6184;
					out<=204;
				end
			end
			297: begin
				if(in == 0) begin
					state<=298;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=4196;
					out<=207;
				end
				if(in == 3) begin
					state<=2296;
					out<=208;
				end
				if(in == 4) begin
					state<=6185;
					out<=209;
				end
			end
			298: begin
				if(in == 0) begin
					state<=299;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=4197;
					out<=212;
				end
				if(in == 3) begin
					state<=2297;
					out<=213;
				end
				if(in == 4) begin
					state<=6186;
					out<=214;
				end
			end
			299: begin
				if(in == 0) begin
					state<=300;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=4198;
					out<=217;
				end
				if(in == 3) begin
					state<=2298;
					out<=218;
				end
				if(in == 4) begin
					state<=6187;
					out<=219;
				end
			end
			300: begin
				if(in == 0) begin
					state<=301;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=4199;
					out<=222;
				end
				if(in == 3) begin
					state<=2299;
					out<=223;
				end
				if(in == 4) begin
					state<=6188;
					out<=224;
				end
			end
			301: begin
				if(in == 0) begin
					state<=302;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=4200;
					out<=227;
				end
				if(in == 3) begin
					state<=2300;
					out<=228;
				end
				if(in == 4) begin
					state<=6189;
					out<=229;
				end
			end
			302: begin
				if(in == 0) begin
					state<=303;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=4201;
					out<=232;
				end
				if(in == 3) begin
					state<=2301;
					out<=233;
				end
				if(in == 4) begin
					state<=6190;
					out<=234;
				end
			end
			303: begin
				if(in == 0) begin
					state<=304;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=4202;
					out<=237;
				end
				if(in == 3) begin
					state<=2302;
					out<=238;
				end
				if(in == 4) begin
					state<=6191;
					out<=239;
				end
			end
			304: begin
				if(in == 0) begin
					state<=305;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=4203;
					out<=242;
				end
				if(in == 3) begin
					state<=2303;
					out<=243;
				end
				if(in == 4) begin
					state<=6192;
					out<=244;
				end
			end
			305: begin
				if(in == 0) begin
					state<=306;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=4204;
					out<=247;
				end
				if(in == 3) begin
					state<=2304;
					out<=248;
				end
				if(in == 4) begin
					state<=6193;
					out<=249;
				end
			end
			306: begin
				if(in == 0) begin
					state<=307;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=4205;
					out<=252;
				end
				if(in == 3) begin
					state<=2305;
					out<=253;
				end
				if(in == 4) begin
					state<=6194;
					out<=254;
				end
			end
			307: begin
				if(in == 0) begin
					state<=308;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=4206;
					out<=1;
				end
				if(in == 3) begin
					state<=2306;
					out<=2;
				end
				if(in == 4) begin
					state<=6195;
					out<=3;
				end
			end
			308: begin
				if(in == 0) begin
					state<=309;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=4207;
					out<=6;
				end
				if(in == 3) begin
					state<=2307;
					out<=7;
				end
				if(in == 4) begin
					state<=6196;
					out<=8;
				end
			end
			309: begin
				if(in == 0) begin
					state<=310;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=4208;
					out<=11;
				end
				if(in == 3) begin
					state<=2308;
					out<=12;
				end
				if(in == 4) begin
					state<=6197;
					out<=13;
				end
			end
			310: begin
				if(in == 0) begin
					state<=311;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=4209;
					out<=16;
				end
				if(in == 3) begin
					state<=2309;
					out<=17;
				end
				if(in == 4) begin
					state<=6198;
					out<=18;
				end
			end
			311: begin
				if(in == 0) begin
					state<=312;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=4210;
					out<=21;
				end
				if(in == 3) begin
					state<=2310;
					out<=22;
				end
				if(in == 4) begin
					state<=6199;
					out<=23;
				end
			end
			312: begin
				if(in == 0) begin
					state<=313;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=4211;
					out<=26;
				end
				if(in == 3) begin
					state<=2311;
					out<=27;
				end
				if(in == 4) begin
					state<=6200;
					out<=28;
				end
			end
			313: begin
				if(in == 0) begin
					state<=314;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=4212;
					out<=31;
				end
				if(in == 3) begin
					state<=2312;
					out<=32;
				end
				if(in == 4) begin
					state<=6201;
					out<=33;
				end
			end
			314: begin
				if(in == 0) begin
					state<=315;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=4213;
					out<=36;
				end
				if(in == 3) begin
					state<=2313;
					out<=37;
				end
				if(in == 4) begin
					state<=6202;
					out<=38;
				end
			end
			315: begin
				if(in == 0) begin
					state<=316;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=4214;
					out<=41;
				end
				if(in == 3) begin
					state<=2314;
					out<=42;
				end
				if(in == 4) begin
					state<=6203;
					out<=43;
				end
			end
			316: begin
				if(in == 0) begin
					state<=317;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=4215;
					out<=46;
				end
				if(in == 3) begin
					state<=2315;
					out<=47;
				end
				if(in == 4) begin
					state<=6204;
					out<=48;
				end
			end
			317: begin
				if(in == 0) begin
					state<=318;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=4216;
					out<=51;
				end
				if(in == 3) begin
					state<=2316;
					out<=52;
				end
				if(in == 4) begin
					state<=6205;
					out<=53;
				end
			end
			318: begin
				if(in == 0) begin
					state<=319;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=4217;
					out<=56;
				end
				if(in == 3) begin
					state<=2317;
					out<=57;
				end
				if(in == 4) begin
					state<=6206;
					out<=58;
				end
			end
			319: begin
				if(in == 0) begin
					state<=320;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=4218;
					out<=61;
				end
				if(in == 3) begin
					state<=2318;
					out<=62;
				end
				if(in == 4) begin
					state<=6207;
					out<=63;
				end
			end
			320: begin
				if(in == 0) begin
					state<=321;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=4219;
					out<=66;
				end
				if(in == 3) begin
					state<=2319;
					out<=67;
				end
				if(in == 4) begin
					state<=6208;
					out<=68;
				end
			end
			321: begin
				if(in == 0) begin
					state<=322;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=4220;
					out<=71;
				end
				if(in == 3) begin
					state<=2320;
					out<=72;
				end
				if(in == 4) begin
					state<=6209;
					out<=73;
				end
			end
			322: begin
				if(in == 0) begin
					state<=323;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=4221;
					out<=76;
				end
				if(in == 3) begin
					state<=2321;
					out<=77;
				end
				if(in == 4) begin
					state<=6210;
					out<=78;
				end
			end
			323: begin
				if(in == 0) begin
					state<=324;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=4222;
					out<=81;
				end
				if(in == 3) begin
					state<=2322;
					out<=82;
				end
				if(in == 4) begin
					state<=6211;
					out<=83;
				end
			end
			324: begin
				if(in == 0) begin
					state<=325;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=4223;
					out<=86;
				end
				if(in == 3) begin
					state<=2323;
					out<=87;
				end
				if(in == 4) begin
					state<=6212;
					out<=88;
				end
			end
			325: begin
				if(in == 0) begin
					state<=326;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=4224;
					out<=91;
				end
				if(in == 3) begin
					state<=2324;
					out<=92;
				end
				if(in == 4) begin
					state<=6213;
					out<=93;
				end
			end
			326: begin
				if(in == 0) begin
					state<=1453;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=5342;
					out<=96;
				end
				if(in == 3) begin
					state<=2898;
					out<=97;
				end
				if(in == 4) begin
					state<=6787;
					out<=98;
				end
			end
			327: begin
				if(in == 0) begin
					state<=328;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=4226;
					out<=101;
				end
				if(in == 3) begin
					state<=2326;
					out<=102;
				end
				if(in == 4) begin
					state<=6215;
					out<=103;
				end
			end
			328: begin
				if(in == 0) begin
					state<=329;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=4227;
					out<=106;
				end
				if(in == 3) begin
					state<=2327;
					out<=107;
				end
				if(in == 4) begin
					state<=6216;
					out<=108;
				end
			end
			329: begin
				if(in == 0) begin
					state<=330;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=4228;
					out<=111;
				end
				if(in == 3) begin
					state<=2328;
					out<=112;
				end
				if(in == 4) begin
					state<=6217;
					out<=113;
				end
			end
			330: begin
				if(in == 0) begin
					state<=331;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=4229;
					out<=116;
				end
				if(in == 3) begin
					state<=2329;
					out<=117;
				end
				if(in == 4) begin
					state<=6218;
					out<=118;
				end
			end
			331: begin
				if(in == 0) begin
					state<=332;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=4230;
					out<=121;
				end
				if(in == 3) begin
					state<=2330;
					out<=122;
				end
				if(in == 4) begin
					state<=6219;
					out<=123;
				end
			end
			332: begin
				if(in == 0) begin
					state<=333;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=4231;
					out<=126;
				end
				if(in == 3) begin
					state<=2331;
					out<=127;
				end
				if(in == 4) begin
					state<=6220;
					out<=128;
				end
			end
			333: begin
				if(in == 0) begin
					state<=334;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=4232;
					out<=131;
				end
				if(in == 3) begin
					state<=2332;
					out<=132;
				end
				if(in == 4) begin
					state<=6221;
					out<=133;
				end
			end
			334: begin
				if(in == 0) begin
					state<=335;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=4233;
					out<=136;
				end
				if(in == 3) begin
					state<=2333;
					out<=137;
				end
				if(in == 4) begin
					state<=6222;
					out<=138;
				end
			end
			335: begin
				if(in == 0) begin
					state<=336;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=4234;
					out<=141;
				end
				if(in == 3) begin
					state<=2334;
					out<=142;
				end
				if(in == 4) begin
					state<=6223;
					out<=143;
				end
			end
			336: begin
				if(in == 0) begin
					state<=337;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=4235;
					out<=146;
				end
				if(in == 3) begin
					state<=2335;
					out<=147;
				end
				if(in == 4) begin
					state<=6224;
					out<=148;
				end
			end
			337: begin
				if(in == 0) begin
					state<=338;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=4236;
					out<=151;
				end
				if(in == 3) begin
					state<=2336;
					out<=152;
				end
				if(in == 4) begin
					state<=6225;
					out<=153;
				end
			end
			338: begin
				if(in == 0) begin
					state<=339;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=4237;
					out<=156;
				end
				if(in == 3) begin
					state<=2337;
					out<=157;
				end
				if(in == 4) begin
					state<=6226;
					out<=158;
				end
			end
			339: begin
				if(in == 0) begin
					state<=340;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=4238;
					out<=161;
				end
				if(in == 3) begin
					state<=2338;
					out<=162;
				end
				if(in == 4) begin
					state<=6227;
					out<=163;
				end
			end
			340: begin
				if(in == 0) begin
					state<=341;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=4239;
					out<=166;
				end
				if(in == 3) begin
					state<=2339;
					out<=167;
				end
				if(in == 4) begin
					state<=6228;
					out<=168;
				end
			end
			341: begin
				if(in == 0) begin
					state<=342;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=4240;
					out<=171;
				end
				if(in == 3) begin
					state<=2340;
					out<=172;
				end
				if(in == 4) begin
					state<=6229;
					out<=173;
				end
			end
			342: begin
				if(in == 0) begin
					state<=343;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=4241;
					out<=176;
				end
				if(in == 3) begin
					state<=2341;
					out<=177;
				end
				if(in == 4) begin
					state<=6230;
					out<=178;
				end
			end
			343: begin
				if(in == 0) begin
					state<=344;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=4242;
					out<=181;
				end
				if(in == 3) begin
					state<=2342;
					out<=182;
				end
				if(in == 4) begin
					state<=6231;
					out<=183;
				end
			end
			344: begin
				if(in == 0) begin
					state<=345;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=4243;
					out<=186;
				end
				if(in == 3) begin
					state<=2343;
					out<=187;
				end
				if(in == 4) begin
					state<=6232;
					out<=188;
				end
			end
			345: begin
				if(in == 0) begin
					state<=346;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=4244;
					out<=191;
				end
				if(in == 3) begin
					state<=2344;
					out<=192;
				end
				if(in == 4) begin
					state<=6233;
					out<=193;
				end
			end
			346: begin
				if(in == 0) begin
					state<=347;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=4245;
					out<=196;
				end
				if(in == 3) begin
					state<=2930;
					out<=197;
				end
				if(in == 4) begin
					state<=6819;
					out<=198;
				end
			end
			347: begin
				if(in == 0) begin
					state<=348;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=4246;
					out<=201;
				end
				if(in == 3) begin
					state<=2931;
					out<=202;
				end
				if(in == 4) begin
					state<=6820;
					out<=203;
				end
			end
			348: begin
				if(in == 0) begin
					state<=349;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=4247;
					out<=206;
				end
				if(in == 3) begin
					state<=2932;
					out<=207;
				end
				if(in == 4) begin
					state<=6821;
					out<=208;
				end
			end
			349: begin
				if(in == 0) begin
					state<=350;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=4248;
					out<=211;
				end
				if(in == 3) begin
					state<=2933;
					out<=212;
				end
				if(in == 4) begin
					state<=6822;
					out<=213;
				end
			end
			350: begin
				if(in == 0) begin
					state<=351;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=4249;
					out<=216;
				end
				if(in == 3) begin
					state<=2934;
					out<=217;
				end
				if(in == 4) begin
					state<=6823;
					out<=218;
				end
			end
			351: begin
				if(in == 0) begin
					state<=352;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=4250;
					out<=221;
				end
				if(in == 3) begin
					state<=2935;
					out<=222;
				end
				if(in == 4) begin
					state<=6824;
					out<=223;
				end
			end
			352: begin
				if(in == 0) begin
					state<=353;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=4251;
					out<=226;
				end
				if(in == 3) begin
					state<=2936;
					out<=227;
				end
				if(in == 4) begin
					state<=6825;
					out<=228;
				end
			end
			353: begin
				if(in == 0) begin
					state<=354;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=4252;
					out<=231;
				end
				if(in == 3) begin
					state<=2937;
					out<=232;
				end
				if(in == 4) begin
					state<=6826;
					out<=233;
				end
			end
			354: begin
				if(in == 0) begin
					state<=355;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=4253;
					out<=236;
				end
				if(in == 3) begin
					state<=2938;
					out<=237;
				end
				if(in == 4) begin
					state<=6827;
					out<=238;
				end
			end
			355: begin
				if(in == 0) begin
					state<=356;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=4254;
					out<=241;
				end
				if(in == 3) begin
					state<=2939;
					out<=242;
				end
				if(in == 4) begin
					state<=6828;
					out<=243;
				end
			end
			356: begin
				if(in == 0) begin
					state<=357;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=4255;
					out<=246;
				end
				if(in == 3) begin
					state<=2940;
					out<=247;
				end
				if(in == 4) begin
					state<=6829;
					out<=248;
				end
			end
			357: begin
				if(in == 0) begin
					state<=358;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=4256;
					out<=251;
				end
				if(in == 3) begin
					state<=2941;
					out<=252;
				end
				if(in == 4) begin
					state<=6830;
					out<=253;
				end
			end
			358: begin
				if(in == 0) begin
					state<=359;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=4257;
					out<=0;
				end
				if(in == 3) begin
					state<=2942;
					out<=1;
				end
				if(in == 4) begin
					state<=6831;
					out<=2;
				end
			end
			359: begin
				if(in == 0) begin
					state<=360;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=4258;
					out<=5;
				end
				if(in == 3) begin
					state<=2943;
					out<=6;
				end
				if(in == 4) begin
					state<=6832;
					out<=7;
				end
			end
			360: begin
				if(in == 0) begin
					state<=361;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=4259;
					out<=10;
				end
				if(in == 3) begin
					state<=2944;
					out<=11;
				end
				if(in == 4) begin
					state<=6833;
					out<=12;
				end
			end
			361: begin
				if(in == 0) begin
					state<=362;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=4260;
					out<=15;
				end
				if(in == 3) begin
					state<=2945;
					out<=16;
				end
				if(in == 4) begin
					state<=6834;
					out<=17;
				end
			end
			362: begin
				if(in == 0) begin
					state<=363;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=4261;
					out<=20;
				end
				if(in == 3) begin
					state<=2946;
					out<=21;
				end
				if(in == 4) begin
					state<=6835;
					out<=22;
				end
			end
			363: begin
				if(in == 0) begin
					state<=364;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=4262;
					out<=25;
				end
				if(in == 3) begin
					state<=2947;
					out<=26;
				end
				if(in == 4) begin
					state<=6836;
					out<=27;
				end
			end
			364: begin
				if(in == 0) begin
					state<=365;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=4263;
					out<=30;
				end
				if(in == 3) begin
					state<=2948;
					out<=31;
				end
				if(in == 4) begin
					state<=6837;
					out<=32;
				end
			end
			365: begin
				if(in == 0) begin
					state<=366;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=4264;
					out<=35;
				end
				if(in == 3) begin
					state<=2949;
					out<=36;
				end
				if(in == 4) begin
					state<=6838;
					out<=37;
				end
			end
			366: begin
				if(in == 0) begin
					state<=367;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=4265;
					out<=40;
				end
				if(in == 3) begin
					state<=2950;
					out<=41;
				end
				if(in == 4) begin
					state<=6839;
					out<=42;
				end
			end
			367: begin
				if(in == 0) begin
					state<=368;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=4266;
					out<=45;
				end
				if(in == 3) begin
					state<=2951;
					out<=46;
				end
				if(in == 4) begin
					state<=6840;
					out<=47;
				end
			end
			368: begin
				if(in == 0) begin
					state<=369;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=4267;
					out<=50;
				end
				if(in == 3) begin
					state<=2952;
					out<=51;
				end
				if(in == 4) begin
					state<=6841;
					out<=52;
				end
			end
			369: begin
				if(in == 0) begin
					state<=370;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=4268;
					out<=55;
				end
				if(in == 3) begin
					state<=2953;
					out<=56;
				end
				if(in == 4) begin
					state<=6842;
					out<=57;
				end
			end
			370: begin
				if(in == 0) begin
					state<=371;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=4269;
					out<=60;
				end
				if(in == 3) begin
					state<=2954;
					out<=61;
				end
				if(in == 4) begin
					state<=6843;
					out<=62;
				end
			end
			371: begin
				if(in == 0) begin
					state<=372;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=4270;
					out<=65;
				end
				if(in == 3) begin
					state<=2955;
					out<=66;
				end
				if(in == 4) begin
					state<=6844;
					out<=67;
				end
			end
			372: begin
				if(in == 0) begin
					state<=373;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=4271;
					out<=70;
				end
				if(in == 3) begin
					state<=2956;
					out<=71;
				end
				if(in == 4) begin
					state<=6845;
					out<=72;
				end
			end
			373: begin
				if(in == 0) begin
					state<=374;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=4272;
					out<=75;
				end
				if(in == 3) begin
					state<=2957;
					out<=76;
				end
				if(in == 4) begin
					state<=6846;
					out<=77;
				end
			end
			374: begin
				if(in == 0) begin
					state<=375;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=4273;
					out<=80;
				end
				if(in == 3) begin
					state<=2958;
					out<=81;
				end
				if(in == 4) begin
					state<=6847;
					out<=82;
				end
			end
			375: begin
				if(in == 0) begin
					state<=376;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=4274;
					out<=85;
				end
				if(in == 3) begin
					state<=2959;
					out<=86;
				end
				if(in == 4) begin
					state<=6848;
					out<=87;
				end
			end
			376: begin
				if(in == 0) begin
					state<=377;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=4275;
					out<=90;
				end
				if(in == 3) begin
					state<=2960;
					out<=91;
				end
				if(in == 4) begin
					state<=6849;
					out<=92;
				end
			end
			377: begin
				if(in == 0) begin
					state<=378;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=4276;
					out<=95;
				end
				if(in == 3) begin
					state<=2961;
					out<=96;
				end
				if(in == 4) begin
					state<=6850;
					out<=97;
				end
			end
			378: begin
				if(in == 0) begin
					state<=379;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=4277;
					out<=100;
				end
				if(in == 3) begin
					state<=2962;
					out<=101;
				end
				if(in == 4) begin
					state<=6851;
					out<=102;
				end
			end
			379: begin
				if(in == 0) begin
					state<=380;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=4278;
					out<=105;
				end
				if(in == 3) begin
					state<=2963;
					out<=106;
				end
				if(in == 4) begin
					state<=6852;
					out<=107;
				end
			end
			380: begin
				if(in == 0) begin
					state<=381;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=4279;
					out<=110;
				end
				if(in == 3) begin
					state<=2964;
					out<=111;
				end
				if(in == 4) begin
					state<=6853;
					out<=112;
				end
			end
			381: begin
				if(in == 0) begin
					state<=382;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=4280;
					out<=115;
				end
				if(in == 3) begin
					state<=2965;
					out<=116;
				end
				if(in == 4) begin
					state<=6854;
					out<=117;
				end
			end
			382: begin
				if(in == 0) begin
					state<=383;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=4281;
					out<=120;
				end
				if(in == 3) begin
					state<=2966;
					out<=121;
				end
				if(in == 4) begin
					state<=6855;
					out<=122;
				end
			end
			383: begin
				if(in == 0) begin
					state<=384;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=4282;
					out<=125;
				end
				if(in == 3) begin
					state<=2967;
					out<=126;
				end
				if(in == 4) begin
					state<=6856;
					out<=127;
				end
			end
			384: begin
				if(in == 0) begin
					state<=385;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=4283;
					out<=130;
				end
				if(in == 3) begin
					state<=2968;
					out<=131;
				end
				if(in == 4) begin
					state<=6857;
					out<=132;
				end
			end
			385: begin
				if(in == 0) begin
					state<=386;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=4284;
					out<=135;
				end
				if(in == 3) begin
					state<=2969;
					out<=136;
				end
				if(in == 4) begin
					state<=6858;
					out<=137;
				end
			end
			386: begin
				if(in == 0) begin
					state<=387;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=4285;
					out<=140;
				end
				if(in == 3) begin
					state<=2970;
					out<=141;
				end
				if(in == 4) begin
					state<=6859;
					out<=142;
				end
			end
			387: begin
				if(in == 0) begin
					state<=388;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=4286;
					out<=145;
				end
				if(in == 3) begin
					state<=2971;
					out<=146;
				end
				if(in == 4) begin
					state<=6860;
					out<=147;
				end
			end
			388: begin
				if(in == 0) begin
					state<=389;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=4287;
					out<=150;
				end
				if(in == 3) begin
					state<=2972;
					out<=151;
				end
				if(in == 4) begin
					state<=6861;
					out<=152;
				end
			end
			389: begin
				if(in == 0) begin
					state<=390;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=4288;
					out<=155;
				end
				if(in == 3) begin
					state<=2973;
					out<=156;
				end
				if(in == 4) begin
					state<=6862;
					out<=157;
				end
			end
			390: begin
				if(in == 0) begin
					state<=391;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=4289;
					out<=160;
				end
				if(in == 3) begin
					state<=2974;
					out<=161;
				end
				if(in == 4) begin
					state<=6863;
					out<=162;
				end
			end
			391: begin
				if(in == 0) begin
					state<=392;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=4290;
					out<=165;
				end
				if(in == 3) begin
					state<=2975;
					out<=166;
				end
				if(in == 4) begin
					state<=6864;
					out<=167;
				end
			end
			392: begin
				if(in == 0) begin
					state<=393;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=4291;
					out<=170;
				end
				if(in == 3) begin
					state<=2976;
					out<=171;
				end
				if(in == 4) begin
					state<=6865;
					out<=172;
				end
			end
			393: begin
				if(in == 0) begin
					state<=394;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=4292;
					out<=175;
				end
				if(in == 3) begin
					state<=2977;
					out<=176;
				end
				if(in == 4) begin
					state<=6866;
					out<=177;
				end
			end
			394: begin
				if(in == 0) begin
					state<=395;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=4293;
					out<=180;
				end
				if(in == 3) begin
					state<=2978;
					out<=181;
				end
				if(in == 4) begin
					state<=6867;
					out<=182;
				end
			end
			395: begin
				if(in == 0) begin
					state<=999;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=4897;
					out<=185;
				end
				if(in == 3) begin
					state<=2979;
					out<=186;
				end
				if(in == 4) begin
					state<=6868;
					out<=187;
				end
			end
			396: begin
				if(in == 0) begin
					state<=397;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=4295;
					out<=190;
				end
				if(in == 3) begin
					state<=3011;
					out<=191;
				end
				if(in == 4) begin
					state<=6900;
					out<=192;
				end
			end
			397: begin
				if(in == 0) begin
					state<=398;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=4296;
					out<=195;
				end
				if(in == 3) begin
					state<=3012;
					out<=196;
				end
				if(in == 4) begin
					state<=6901;
					out<=197;
				end
			end
			398: begin
				if(in == 0) begin
					state<=399;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=4297;
					out<=200;
				end
				if(in == 3) begin
					state<=3013;
					out<=201;
				end
				if(in == 4) begin
					state<=6902;
					out<=202;
				end
			end
			399: begin
				if(in == 0) begin
					state<=400;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=4298;
					out<=205;
				end
				if(in == 3) begin
					state<=3014;
					out<=206;
				end
				if(in == 4) begin
					state<=6903;
					out<=207;
				end
			end
			400: begin
				if(in == 0) begin
					state<=401;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=4299;
					out<=210;
				end
				if(in == 3) begin
					state<=3015;
					out<=211;
				end
				if(in == 4) begin
					state<=6904;
					out<=212;
				end
			end
			401: begin
				if(in == 0) begin
					state<=402;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=4300;
					out<=215;
				end
				if(in == 3) begin
					state<=3016;
					out<=216;
				end
				if(in == 4) begin
					state<=6905;
					out<=217;
				end
			end
			402: begin
				if(in == 0) begin
					state<=403;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=4301;
					out<=220;
				end
				if(in == 3) begin
					state<=3017;
					out<=221;
				end
				if(in == 4) begin
					state<=6906;
					out<=222;
				end
			end
			403: begin
				if(in == 0) begin
					state<=404;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=4302;
					out<=225;
				end
				if(in == 3) begin
					state<=3018;
					out<=226;
				end
				if(in == 4) begin
					state<=6907;
					out<=227;
				end
			end
			404: begin
				if(in == 0) begin
					state<=405;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=4303;
					out<=230;
				end
				if(in == 3) begin
					state<=3019;
					out<=231;
				end
				if(in == 4) begin
					state<=6908;
					out<=232;
				end
			end
			405: begin
				if(in == 0) begin
					state<=406;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=4304;
					out<=235;
				end
				if(in == 3) begin
					state<=3020;
					out<=236;
				end
				if(in == 4) begin
					state<=6909;
					out<=237;
				end
			end
			406: begin
				if(in == 0) begin
					state<=407;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=4305;
					out<=240;
				end
				if(in == 3) begin
					state<=3021;
					out<=241;
				end
				if(in == 4) begin
					state<=6910;
					out<=242;
				end
			end
			407: begin
				if(in == 0) begin
					state<=408;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=4306;
					out<=245;
				end
				if(in == 3) begin
					state<=3022;
					out<=246;
				end
				if(in == 4) begin
					state<=6911;
					out<=247;
				end
			end
			408: begin
				if(in == 0) begin
					state<=409;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=4307;
					out<=250;
				end
				if(in == 3) begin
					state<=3023;
					out<=251;
				end
				if(in == 4) begin
					state<=6912;
					out<=252;
				end
			end
			409: begin
				if(in == 0) begin
					state<=410;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=4308;
					out<=255;
				end
				if(in == 3) begin
					state<=3024;
					out<=0;
				end
				if(in == 4) begin
					state<=6913;
					out<=1;
				end
			end
			410: begin
				if(in == 0) begin
					state<=411;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=4309;
					out<=4;
				end
				if(in == 3) begin
					state<=3025;
					out<=5;
				end
				if(in == 4) begin
					state<=6914;
					out<=6;
				end
			end
			411: begin
				if(in == 0) begin
					state<=412;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=4310;
					out<=9;
				end
				if(in == 3) begin
					state<=3026;
					out<=10;
				end
				if(in == 4) begin
					state<=6915;
					out<=11;
				end
			end
			412: begin
				if(in == 0) begin
					state<=413;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=4311;
					out<=14;
				end
				if(in == 3) begin
					state<=3027;
					out<=15;
				end
				if(in == 4) begin
					state<=6916;
					out<=16;
				end
			end
			413: begin
				if(in == 0) begin
					state<=414;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=4312;
					out<=19;
				end
				if(in == 3) begin
					state<=3028;
					out<=20;
				end
				if(in == 4) begin
					state<=6917;
					out<=21;
				end
			end
			414: begin
				if(in == 0) begin
					state<=1030;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=4928;
					out<=24;
				end
				if(in == 3) begin
					state<=3029;
					out<=25;
				end
				if(in == 4) begin
					state<=6918;
					out<=26;
				end
			end
			415: begin
				if(in == 0) begin
					state<=416;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=4314;
					out<=29;
				end
				if(in == 3) begin
					state<=2414;
					out<=30;
				end
				if(in == 4) begin
					state<=6303;
					out<=31;
				end
			end
			416: begin
				if(in == 0) begin
					state<=417;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=4315;
					out<=34;
				end
				if(in == 3) begin
					state<=2415;
					out<=35;
				end
				if(in == 4) begin
					state<=6304;
					out<=36;
				end
			end
			417: begin
				if(in == 0) begin
					state<=418;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=4316;
					out<=39;
				end
				if(in == 3) begin
					state<=2416;
					out<=40;
				end
				if(in == 4) begin
					state<=6305;
					out<=41;
				end
			end
			418: begin
				if(in == 0) begin
					state<=419;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=4317;
					out<=44;
				end
				if(in == 3) begin
					state<=2417;
					out<=45;
				end
				if(in == 4) begin
					state<=6306;
					out<=46;
				end
			end
			419: begin
				if(in == 0) begin
					state<=420;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=4318;
					out<=49;
				end
				if(in == 3) begin
					state<=2418;
					out<=50;
				end
				if(in == 4) begin
					state<=6307;
					out<=51;
				end
			end
			420: begin
				if(in == 0) begin
					state<=421;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=4319;
					out<=54;
				end
				if(in == 3) begin
					state<=2419;
					out<=55;
				end
				if(in == 4) begin
					state<=6308;
					out<=56;
				end
			end
			421: begin
				if(in == 0) begin
					state<=422;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=4320;
					out<=59;
				end
				if(in == 3) begin
					state<=2420;
					out<=60;
				end
				if(in == 4) begin
					state<=6309;
					out<=61;
				end
			end
			422: begin
				if(in == 0) begin
					state<=423;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=4321;
					out<=64;
				end
				if(in == 3) begin
					state<=2421;
					out<=65;
				end
				if(in == 4) begin
					state<=6310;
					out<=66;
				end
			end
			423: begin
				if(in == 0) begin
					state<=424;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=4322;
					out<=69;
				end
				if(in == 3) begin
					state<=2422;
					out<=70;
				end
				if(in == 4) begin
					state<=6311;
					out<=71;
				end
			end
			424: begin
				if(in == 0) begin
					state<=425;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=4323;
					out<=74;
				end
				if(in == 3) begin
					state<=2423;
					out<=75;
				end
				if(in == 4) begin
					state<=6312;
					out<=76;
				end
			end
			425: begin
				if(in == 0) begin
					state<=426;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=4324;
					out<=79;
				end
				if(in == 3) begin
					state<=2424;
					out<=80;
				end
				if(in == 4) begin
					state<=6313;
					out<=81;
				end
			end
			426: begin
				if(in == 0) begin
					state<=427;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=4325;
					out<=84;
				end
				if(in == 3) begin
					state<=2425;
					out<=85;
				end
				if(in == 4) begin
					state<=6314;
					out<=86;
				end
			end
			427: begin
				if(in == 0) begin
					state<=428;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=4326;
					out<=89;
				end
				if(in == 3) begin
					state<=2426;
					out<=90;
				end
				if(in == 4) begin
					state<=6315;
					out<=91;
				end
			end
			428: begin
				if(in == 0) begin
					state<=429;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=4327;
					out<=94;
				end
				if(in == 3) begin
					state<=2427;
					out<=95;
				end
				if(in == 4) begin
					state<=6316;
					out<=96;
				end
			end
			429: begin
				if(in == 0) begin
					state<=430;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=4328;
					out<=99;
				end
				if(in == 3) begin
					state<=2428;
					out<=100;
				end
				if(in == 4) begin
					state<=6317;
					out<=101;
				end
			end
			430: begin
				if(in == 0) begin
					state<=431;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=4329;
					out<=104;
				end
				if(in == 3) begin
					state<=2429;
					out<=105;
				end
				if(in == 4) begin
					state<=6318;
					out<=106;
				end
			end
			431: begin
				if(in == 0) begin
					state<=432;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=4330;
					out<=109;
				end
				if(in == 3) begin
					state<=2430;
					out<=110;
				end
				if(in == 4) begin
					state<=6319;
					out<=111;
				end
			end
			432: begin
				if(in == 0) begin
					state<=433;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=4331;
					out<=114;
				end
				if(in == 3) begin
					state<=2431;
					out<=115;
				end
				if(in == 4) begin
					state<=6320;
					out<=116;
				end
			end
			433: begin
				if(in == 0) begin
					state<=434;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=4332;
					out<=119;
				end
				if(in == 3) begin
					state<=2432;
					out<=120;
				end
				if(in == 4) begin
					state<=6321;
					out<=121;
				end
			end
			434: begin
				if(in == 0) begin
					state<=435;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=4333;
					out<=124;
				end
				if(in == 3) begin
					state<=2433;
					out<=125;
				end
				if(in == 4) begin
					state<=6322;
					out<=126;
				end
			end
			435: begin
				if(in == 0) begin
					state<=436;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=4334;
					out<=129;
				end
				if(in == 3) begin
					state<=2434;
					out<=130;
				end
				if(in == 4) begin
					state<=6323;
					out<=131;
				end
			end
			436: begin
				if(in == 0) begin
					state<=437;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=4335;
					out<=134;
				end
				if(in == 3) begin
					state<=2435;
					out<=135;
				end
				if(in == 4) begin
					state<=6324;
					out<=136;
				end
			end
			437: begin
				if(in == 0) begin
					state<=438;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=4336;
					out<=139;
				end
				if(in == 3) begin
					state<=2436;
					out<=140;
				end
				if(in == 4) begin
					state<=6325;
					out<=141;
				end
			end
			438: begin
				if(in == 0) begin
					state<=439;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=4337;
					out<=144;
				end
				if(in == 3) begin
					state<=2437;
					out<=145;
				end
				if(in == 4) begin
					state<=6326;
					out<=146;
				end
			end
			439: begin
				if(in == 0) begin
					state<=440;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=4338;
					out<=149;
				end
				if(in == 3) begin
					state<=2438;
					out<=150;
				end
				if(in == 4) begin
					state<=6327;
					out<=151;
				end
			end
			440: begin
				if(in == 0) begin
					state<=441;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=4339;
					out<=154;
				end
				if(in == 3) begin
					state<=2439;
					out<=155;
				end
				if(in == 4) begin
					state<=6328;
					out<=156;
				end
			end
			441: begin
				if(in == 0) begin
					state<=442;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=4340;
					out<=159;
				end
				if(in == 3) begin
					state<=2440;
					out<=160;
				end
				if(in == 4) begin
					state<=6329;
					out<=161;
				end
			end
			442: begin
				if(in == 0) begin
					state<=443;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=4341;
					out<=164;
				end
				if(in == 3) begin
					state<=2441;
					out<=165;
				end
				if(in == 4) begin
					state<=6330;
					out<=166;
				end
			end
			443: begin
				if(in == 0) begin
					state<=444;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=4342;
					out<=169;
				end
				if(in == 3) begin
					state<=2442;
					out<=170;
				end
				if(in == 4) begin
					state<=6331;
					out<=171;
				end
			end
			444: begin
				if(in == 0) begin
					state<=445;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=4343;
					out<=174;
				end
				if(in == 3) begin
					state<=2443;
					out<=175;
				end
				if(in == 4) begin
					state<=6332;
					out<=176;
				end
			end
			445: begin
				if(in == 0) begin
					state<=446;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=4344;
					out<=179;
				end
				if(in == 3) begin
					state<=2444;
					out<=180;
				end
				if(in == 4) begin
					state<=6333;
					out<=181;
				end
			end
			446: begin
				if(in == 0) begin
					state<=447;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=4345;
					out<=184;
				end
				if(in == 3) begin
					state<=2445;
					out<=185;
				end
				if(in == 4) begin
					state<=6334;
					out<=186;
				end
			end
			447: begin
				if(in == 0) begin
					state<=448;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=4346;
					out<=189;
				end
				if(in == 3) begin
					state<=2446;
					out<=190;
				end
				if(in == 4) begin
					state<=6335;
					out<=191;
				end
			end
			448: begin
				if(in == 0) begin
					state<=449;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=4347;
					out<=194;
				end
				if(in == 3) begin
					state<=2447;
					out<=195;
				end
				if(in == 4) begin
					state<=6336;
					out<=196;
				end
			end
			449: begin
				if(in == 0) begin
					state<=450;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=4348;
					out<=199;
				end
				if(in == 3) begin
					state<=2448;
					out<=200;
				end
				if(in == 4) begin
					state<=6337;
					out<=201;
				end
			end
			450: begin
				if(in == 0) begin
					state<=451;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=4349;
					out<=204;
				end
				if(in == 3) begin
					state<=2449;
					out<=205;
				end
				if(in == 4) begin
					state<=6338;
					out<=206;
				end
			end
			451: begin
				if(in == 0) begin
					state<=452;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=4350;
					out<=209;
				end
				if(in == 3) begin
					state<=2450;
					out<=210;
				end
				if(in == 4) begin
					state<=6339;
					out<=211;
				end
			end
			452: begin
				if(in == 0) begin
					state<=453;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=4351;
					out<=214;
				end
				if(in == 3) begin
					state<=2451;
					out<=215;
				end
				if(in == 4) begin
					state<=6340;
					out<=216;
				end
			end
			453: begin
				if(in == 0) begin
					state<=454;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=4352;
					out<=219;
				end
				if(in == 3) begin
					state<=2452;
					out<=220;
				end
				if(in == 4) begin
					state<=6341;
					out<=221;
				end
			end
			454: begin
				if(in == 0) begin
					state<=455;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=4353;
					out<=224;
				end
				if(in == 3) begin
					state<=2453;
					out<=225;
				end
				if(in == 4) begin
					state<=6342;
					out<=226;
				end
			end
			455: begin
				if(in == 0) begin
					state<=456;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=4354;
					out<=229;
				end
				if(in == 3) begin
					state<=2454;
					out<=230;
				end
				if(in == 4) begin
					state<=6343;
					out<=231;
				end
			end
			456: begin
				if(in == 0) begin
					state<=457;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=4355;
					out<=234;
				end
				if(in == 3) begin
					state<=2455;
					out<=235;
				end
				if(in == 4) begin
					state<=6344;
					out<=236;
				end
			end
			457: begin
				if(in == 0) begin
					state<=458;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=4356;
					out<=239;
				end
				if(in == 3) begin
					state<=2456;
					out<=240;
				end
				if(in == 4) begin
					state<=6345;
					out<=241;
				end
			end
			458: begin
				if(in == 0) begin
					state<=459;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=4357;
					out<=244;
				end
				if(in == 3) begin
					state<=2457;
					out<=245;
				end
				if(in == 4) begin
					state<=6346;
					out<=246;
				end
			end
			459: begin
				if(in == 0) begin
					state<=460;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=4358;
					out<=249;
				end
				if(in == 3) begin
					state<=2458;
					out<=250;
				end
				if(in == 4) begin
					state<=6347;
					out<=251;
				end
			end
			460: begin
				if(in == 0) begin
					state<=461;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=4359;
					out<=254;
				end
				if(in == 3) begin
					state<=2459;
					out<=255;
				end
				if(in == 4) begin
					state<=6348;
					out<=0;
				end
			end
			461: begin
				if(in == 0) begin
					state<=462;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=4360;
					out<=3;
				end
				if(in == 3) begin
					state<=2460;
					out<=4;
				end
				if(in == 4) begin
					state<=6349;
					out<=5;
				end
			end
			462: begin
				if(in == 0) begin
					state<=463;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=4361;
					out<=8;
				end
				if(in == 3) begin
					state<=2461;
					out<=9;
				end
				if(in == 4) begin
					state<=6350;
					out<=10;
				end
			end
			463: begin
				if(in == 0) begin
					state<=464;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=4362;
					out<=13;
				end
				if(in == 3) begin
					state<=2462;
					out<=14;
				end
				if(in == 4) begin
					state<=6351;
					out<=15;
				end
			end
			464: begin
				if(in == 0) begin
					state<=1484;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=5373;
					out<=18;
				end
				if(in == 3) begin
					state<=3416;
					out<=19;
				end
				if(in == 4) begin
					state<=7305;
					out<=20;
				end
			end
			465: begin
				if(in == 0) begin
					state<=466;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=4364;
					out<=23;
				end
				if(in == 3) begin
					state<=2464;
					out<=24;
				end
				if(in == 4) begin
					state<=6353;
					out<=25;
				end
			end
			466: begin
				if(in == 0) begin
					state<=467;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=4365;
					out<=28;
				end
				if(in == 3) begin
					state<=2465;
					out<=29;
				end
				if(in == 4) begin
					state<=6354;
					out<=30;
				end
			end
			467: begin
				if(in == 0) begin
					state<=468;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=4366;
					out<=33;
				end
				if(in == 3) begin
					state<=2466;
					out<=34;
				end
				if(in == 4) begin
					state<=6355;
					out<=35;
				end
			end
			468: begin
				if(in == 0) begin
					state<=469;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=4367;
					out<=38;
				end
				if(in == 3) begin
					state<=2467;
					out<=39;
				end
				if(in == 4) begin
					state<=6356;
					out<=40;
				end
			end
			469: begin
				if(in == 0) begin
					state<=470;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=4368;
					out<=43;
				end
				if(in == 3) begin
					state<=2468;
					out<=44;
				end
				if(in == 4) begin
					state<=6357;
					out<=45;
				end
			end
			470: begin
				if(in == 0) begin
					state<=471;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=4369;
					out<=48;
				end
				if(in == 3) begin
					state<=2469;
					out<=49;
				end
				if(in == 4) begin
					state<=6358;
					out<=50;
				end
			end
			471: begin
				if(in == 0) begin
					state<=472;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=4370;
					out<=53;
				end
				if(in == 3) begin
					state<=2470;
					out<=54;
				end
				if(in == 4) begin
					state<=6359;
					out<=55;
				end
			end
			472: begin
				if(in == 0) begin
					state<=473;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=4371;
					out<=58;
				end
				if(in == 3) begin
					state<=2471;
					out<=59;
				end
				if(in == 4) begin
					state<=6360;
					out<=60;
				end
			end
			473: begin
				if(in == 0) begin
					state<=474;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=4372;
					out<=63;
				end
				if(in == 3) begin
					state<=2472;
					out<=64;
				end
				if(in == 4) begin
					state<=6361;
					out<=65;
				end
			end
			474: begin
				if(in == 0) begin
					state<=475;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=4373;
					out<=68;
				end
				if(in == 3) begin
					state<=2473;
					out<=69;
				end
				if(in == 4) begin
					state<=6362;
					out<=70;
				end
			end
			475: begin
				if(in == 0) begin
					state<=476;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=4374;
					out<=73;
				end
				if(in == 3) begin
					state<=2474;
					out<=74;
				end
				if(in == 4) begin
					state<=6363;
					out<=75;
				end
			end
			476: begin
				if(in == 0) begin
					state<=477;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=4375;
					out<=78;
				end
				if(in == 3) begin
					state<=2475;
					out<=79;
				end
				if(in == 4) begin
					state<=6364;
					out<=80;
				end
			end
			477: begin
				if(in == 0) begin
					state<=478;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=4376;
					out<=83;
				end
				if(in == 3) begin
					state<=2476;
					out<=84;
				end
				if(in == 4) begin
					state<=6365;
					out<=85;
				end
			end
			478: begin
				if(in == 0) begin
					state<=479;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=4377;
					out<=88;
				end
				if(in == 3) begin
					state<=2477;
					out<=89;
				end
				if(in == 4) begin
					state<=6366;
					out<=90;
				end
			end
			479: begin
				if(in == 0) begin
					state<=480;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=4378;
					out<=93;
				end
				if(in == 3) begin
					state<=2478;
					out<=94;
				end
				if(in == 4) begin
					state<=6367;
					out<=95;
				end
			end
			480: begin
				if(in == 0) begin
					state<=481;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=4379;
					out<=98;
				end
				if(in == 3) begin
					state<=2479;
					out<=99;
				end
				if(in == 4) begin
					state<=6368;
					out<=100;
				end
			end
			481: begin
				if(in == 0) begin
					state<=482;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=4380;
					out<=103;
				end
				if(in == 3) begin
					state<=2480;
					out<=104;
				end
				if(in == 4) begin
					state<=6369;
					out<=105;
				end
			end
			482: begin
				if(in == 0) begin
					state<=483;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=4381;
					out<=108;
				end
				if(in == 3) begin
					state<=2481;
					out<=109;
				end
				if(in == 4) begin
					state<=6370;
					out<=110;
				end
			end
			483: begin
				if(in == 0) begin
					state<=484;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=4382;
					out<=113;
				end
				if(in == 3) begin
					state<=2482;
					out<=114;
				end
				if(in == 4) begin
					state<=6371;
					out<=115;
				end
			end
			484: begin
				if(in == 0) begin
					state<=485;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=4383;
					out<=118;
				end
				if(in == 3) begin
					state<=2483;
					out<=119;
				end
				if(in == 4) begin
					state<=6372;
					out<=120;
				end
			end
			485: begin
				if(in == 0) begin
					state<=486;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=4384;
					out<=123;
				end
				if(in == 3) begin
					state<=2484;
					out<=124;
				end
				if(in == 4) begin
					state<=6373;
					out<=125;
				end
			end
			486: begin
				if(in == 0) begin
					state<=487;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=4385;
					out<=128;
				end
				if(in == 3) begin
					state<=2485;
					out<=129;
				end
				if(in == 4) begin
					state<=6374;
					out<=130;
				end
			end
			487: begin
				if(in == 0) begin
					state<=488;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=4386;
					out<=133;
				end
				if(in == 3) begin
					state<=2486;
					out<=134;
				end
				if(in == 4) begin
					state<=6375;
					out<=135;
				end
			end
			488: begin
				if(in == 0) begin
					state<=489;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=4387;
					out<=138;
				end
				if(in == 3) begin
					state<=2487;
					out<=139;
				end
				if(in == 4) begin
					state<=6376;
					out<=140;
				end
			end
			489: begin
				if(in == 0) begin
					state<=490;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=4388;
					out<=143;
				end
				if(in == 3) begin
					state<=2488;
					out<=144;
				end
				if(in == 4) begin
					state<=6377;
					out<=145;
				end
			end
			490: begin
				if(in == 0) begin
					state<=491;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=4389;
					out<=148;
				end
				if(in == 3) begin
					state<=2489;
					out<=149;
				end
				if(in == 4) begin
					state<=6378;
					out<=150;
				end
			end
			491: begin
				if(in == 0) begin
					state<=492;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=4390;
					out<=153;
				end
				if(in == 3) begin
					state<=2490;
					out<=154;
				end
				if(in == 4) begin
					state<=6379;
					out<=155;
				end
			end
			492: begin
				if(in == 0) begin
					state<=493;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=4391;
					out<=158;
				end
				if(in == 3) begin
					state<=2491;
					out<=159;
				end
				if(in == 4) begin
					state<=6380;
					out<=160;
				end
			end
			493: begin
				if(in == 0) begin
					state<=494;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=4392;
					out<=163;
				end
				if(in == 3) begin
					state<=2492;
					out<=164;
				end
				if(in == 4) begin
					state<=6381;
					out<=165;
				end
			end
			494: begin
				if(in == 0) begin
					state<=495;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=4393;
					out<=168;
				end
				if(in == 3) begin
					state<=2493;
					out<=169;
				end
				if(in == 4) begin
					state<=6382;
					out<=170;
				end
			end
			495: begin
				if(in == 0) begin
					state<=496;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=4394;
					out<=173;
				end
				if(in == 3) begin
					state<=2494;
					out<=174;
				end
				if(in == 4) begin
					state<=6383;
					out<=175;
				end
			end
			496: begin
				if(in == 0) begin
					state<=497;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=4395;
					out<=178;
				end
				if(in == 3) begin
					state<=2495;
					out<=179;
				end
				if(in == 4) begin
					state<=6384;
					out<=180;
				end
			end
			497: begin
				if(in == 0) begin
					state<=498;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=4396;
					out<=183;
				end
				if(in == 3) begin
					state<=2496;
					out<=184;
				end
				if(in == 4) begin
					state<=6385;
					out<=185;
				end
			end
			498: begin
				if(in == 0) begin
					state<=499;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=4397;
					out<=188;
				end
				if(in == 3) begin
					state<=2497;
					out<=189;
				end
				if(in == 4) begin
					state<=6386;
					out<=190;
				end
			end
			499: begin
				if(in == 0) begin
					state<=500;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=4398;
					out<=193;
				end
				if(in == 3) begin
					state<=2498;
					out<=194;
				end
				if(in == 4) begin
					state<=6387;
					out<=195;
				end
			end
			500: begin
				if(in == 0) begin
					state<=501;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=4399;
					out<=198;
				end
				if(in == 3) begin
					state<=2499;
					out<=199;
				end
				if(in == 4) begin
					state<=6388;
					out<=200;
				end
			end
			501: begin
				if(in == 0) begin
					state<=502;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=4400;
					out<=203;
				end
				if(in == 3) begin
					state<=2500;
					out<=204;
				end
				if(in == 4) begin
					state<=6389;
					out<=205;
				end
			end
			502: begin
				if(in == 0) begin
					state<=503;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=4401;
					out<=208;
				end
				if(in == 3) begin
					state<=2501;
					out<=209;
				end
				if(in == 4) begin
					state<=6390;
					out<=210;
				end
			end
			503: begin
				if(in == 0) begin
					state<=504;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=4402;
					out<=213;
				end
				if(in == 3) begin
					state<=2502;
					out<=214;
				end
				if(in == 4) begin
					state<=6391;
					out<=215;
				end
			end
			504: begin
				if(in == 0) begin
					state<=505;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=4403;
					out<=218;
				end
				if(in == 3) begin
					state<=2503;
					out<=219;
				end
				if(in == 4) begin
					state<=6392;
					out<=220;
				end
			end
			505: begin
				if(in == 0) begin
					state<=506;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=4404;
					out<=223;
				end
				if(in == 3) begin
					state<=2504;
					out<=224;
				end
				if(in == 4) begin
					state<=6393;
					out<=225;
				end
			end
			506: begin
				if(in == 0) begin
					state<=507;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=4405;
					out<=228;
				end
				if(in == 3) begin
					state<=2505;
					out<=229;
				end
				if(in == 4) begin
					state<=6394;
					out<=230;
				end
			end
			507: begin
				if(in == 0) begin
					state<=508;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=4406;
					out<=233;
				end
				if(in == 3) begin
					state<=2506;
					out<=234;
				end
				if(in == 4) begin
					state<=6395;
					out<=235;
				end
			end
			508: begin
				if(in == 0) begin
					state<=509;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=4407;
					out<=238;
				end
				if(in == 3) begin
					state<=2507;
					out<=239;
				end
				if(in == 4) begin
					state<=6396;
					out<=240;
				end
			end
			509: begin
				if(in == 0) begin
					state<=510;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=4408;
					out<=243;
				end
				if(in == 3) begin
					state<=2508;
					out<=244;
				end
				if(in == 4) begin
					state<=6397;
					out<=245;
				end
			end
			510: begin
				if(in == 0) begin
					state<=511;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=4409;
					out<=248;
				end
				if(in == 3) begin
					state<=2509;
					out<=249;
				end
				if(in == 4) begin
					state<=6398;
					out<=250;
				end
			end
			511: begin
				if(in == 0) begin
					state<=512;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=4410;
					out<=253;
				end
				if(in == 3) begin
					state<=2510;
					out<=254;
				end
				if(in == 4) begin
					state<=6399;
					out<=255;
				end
			end
			512: begin
				if(in == 0) begin
					state<=513;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=4411;
					out<=2;
				end
				if(in == 3) begin
					state<=2511;
					out<=3;
				end
				if(in == 4) begin
					state<=6400;
					out<=4;
				end
			end
			513: begin
				if(in == 0) begin
					state<=514;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=4412;
					out<=7;
				end
				if(in == 3) begin
					state<=2512;
					out<=8;
				end
				if(in == 4) begin
					state<=6401;
					out<=9;
				end
			end
			514: begin
				if(in == 0) begin
					state<=515;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=4413;
					out<=12;
				end
				if(in == 3) begin
					state<=2513;
					out<=13;
				end
				if(in == 4) begin
					state<=6402;
					out<=14;
				end
			end
			515: begin
				if(in == 0) begin
					state<=516;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=4414;
					out<=17;
				end
				if(in == 3) begin
					state<=2514;
					out<=18;
				end
				if(in == 4) begin
					state<=6403;
					out<=19;
				end
			end
			516: begin
				if(in == 0) begin
					state<=517;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=4415;
					out<=22;
				end
				if(in == 3) begin
					state<=2515;
					out<=23;
				end
				if(in == 4) begin
					state<=6404;
					out<=24;
				end
			end
			517: begin
				if(in == 0) begin
					state<=518;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=4416;
					out<=27;
				end
				if(in == 3) begin
					state<=2516;
					out<=28;
				end
				if(in == 4) begin
					state<=6405;
					out<=29;
				end
			end
			518: begin
				if(in == 0) begin
					state<=519;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=4417;
					out<=32;
				end
				if(in == 3) begin
					state<=2517;
					out<=33;
				end
				if(in == 4) begin
					state<=6406;
					out<=34;
				end
			end
			519: begin
				if(in == 0) begin
					state<=520;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=4418;
					out<=37;
				end
				if(in == 3) begin
					state<=2518;
					out<=38;
				end
				if(in == 4) begin
					state<=6407;
					out<=39;
				end
			end
			520: begin
				if(in == 0) begin
					state<=521;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=4419;
					out<=42;
				end
				if(in == 3) begin
					state<=2519;
					out<=43;
				end
				if(in == 4) begin
					state<=6408;
					out<=44;
				end
			end
			521: begin
				if(in == 0) begin
					state<=522;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=4420;
					out<=47;
				end
				if(in == 3) begin
					state<=2520;
					out<=48;
				end
				if(in == 4) begin
					state<=6409;
					out<=49;
				end
			end
			522: begin
				if(in == 0) begin
					state<=523;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=4421;
					out<=52;
				end
				if(in == 3) begin
					state<=2521;
					out<=53;
				end
				if(in == 4) begin
					state<=6410;
					out<=54;
				end
			end
			523: begin
				if(in == 0) begin
					state<=524;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=4422;
					out<=57;
				end
				if(in == 3) begin
					state<=2522;
					out<=58;
				end
				if(in == 4) begin
					state<=6411;
					out<=59;
				end
			end
			524: begin
				if(in == 0) begin
					state<=525;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=4423;
					out<=62;
				end
				if(in == 3) begin
					state<=2523;
					out<=63;
				end
				if(in == 4) begin
					state<=6412;
					out<=64;
				end
			end
			525: begin
				if(in == 0) begin
					state<=526;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=4424;
					out<=67;
				end
				if(in == 3) begin
					state<=2524;
					out<=68;
				end
				if(in == 4) begin
					state<=6413;
					out<=69;
				end
			end
			526: begin
				if(in == 0) begin
					state<=527;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=4425;
					out<=72;
				end
				if(in == 3) begin
					state<=2525;
					out<=73;
				end
				if(in == 4) begin
					state<=6414;
					out<=74;
				end
			end
			527: begin
				if(in == 0) begin
					state<=528;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=4426;
					out<=77;
				end
				if(in == 3) begin
					state<=2526;
					out<=78;
				end
				if(in == 4) begin
					state<=6415;
					out<=79;
				end
			end
			528: begin
				if(in == 0) begin
					state<=529;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=4427;
					out<=82;
				end
				if(in == 3) begin
					state<=2527;
					out<=83;
				end
				if(in == 4) begin
					state<=6416;
					out<=84;
				end
			end
			529: begin
				if(in == 0) begin
					state<=530;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=4428;
					out<=87;
				end
				if(in == 3) begin
					state<=2528;
					out<=88;
				end
				if(in == 4) begin
					state<=6417;
					out<=89;
				end
			end
			530: begin
				if(in == 0) begin
					state<=531;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=4429;
					out<=92;
				end
				if(in == 3) begin
					state<=2529;
					out<=93;
				end
				if(in == 4) begin
					state<=6418;
					out<=94;
				end
			end
			531: begin
				if(in == 0) begin
					state<=532;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=4430;
					out<=97;
				end
				if(in == 3) begin
					state<=2530;
					out<=98;
				end
				if(in == 4) begin
					state<=6419;
					out<=99;
				end
			end
			532: begin
				if(in == 0) begin
					state<=533;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=4431;
					out<=102;
				end
				if(in == 3) begin
					state<=2531;
					out<=103;
				end
				if(in == 4) begin
					state<=6420;
					out<=104;
				end
			end
			533: begin
				if(in == 0) begin
					state<=1515;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=5404;
					out<=107;
				end
				if(in == 3) begin
					state<=3447;
					out<=108;
				end
				if(in == 4) begin
					state<=7336;
					out<=109;
				end
			end
			534: begin
				if(in == 0) begin
					state<=535;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=4433;
					out<=112;
				end
				if(in == 3) begin
					state<=2533;
					out<=113;
				end
				if(in == 4) begin
					state<=6422;
					out<=114;
				end
			end
			535: begin
				if(in == 0) begin
					state<=536;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=4434;
					out<=117;
				end
				if(in == 3) begin
					state<=2534;
					out<=118;
				end
				if(in == 4) begin
					state<=6423;
					out<=119;
				end
			end
			536: begin
				if(in == 0) begin
					state<=537;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=4435;
					out<=122;
				end
				if(in == 3) begin
					state<=2535;
					out<=123;
				end
				if(in == 4) begin
					state<=6424;
					out<=124;
				end
			end
			537: begin
				if(in == 0) begin
					state<=538;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=4436;
					out<=127;
				end
				if(in == 3) begin
					state<=2536;
					out<=128;
				end
				if(in == 4) begin
					state<=6425;
					out<=129;
				end
			end
			538: begin
				if(in == 0) begin
					state<=539;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=4437;
					out<=132;
				end
				if(in == 3) begin
					state<=2537;
					out<=133;
				end
				if(in == 4) begin
					state<=6426;
					out<=134;
				end
			end
			539: begin
				if(in == 0) begin
					state<=540;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=4438;
					out<=137;
				end
				if(in == 3) begin
					state<=2538;
					out<=138;
				end
				if(in == 4) begin
					state<=6427;
					out<=139;
				end
			end
			540: begin
				if(in == 0) begin
					state<=541;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=4439;
					out<=142;
				end
				if(in == 3) begin
					state<=2539;
					out<=143;
				end
				if(in == 4) begin
					state<=6428;
					out<=144;
				end
			end
			541: begin
				if(in == 0) begin
					state<=542;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=4440;
					out<=147;
				end
				if(in == 3) begin
					state<=2540;
					out<=148;
				end
				if(in == 4) begin
					state<=6429;
					out<=149;
				end
			end
			542: begin
				if(in == 0) begin
					state<=543;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=4441;
					out<=152;
				end
				if(in == 3) begin
					state<=2541;
					out<=153;
				end
				if(in == 4) begin
					state<=6430;
					out<=154;
				end
			end
			543: begin
				if(in == 0) begin
					state<=544;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=4442;
					out<=157;
				end
				if(in == 3) begin
					state<=2542;
					out<=158;
				end
				if(in == 4) begin
					state<=6431;
					out<=159;
				end
			end
			544: begin
				if(in == 0) begin
					state<=545;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=4443;
					out<=162;
				end
				if(in == 3) begin
					state<=2543;
					out<=163;
				end
				if(in == 4) begin
					state<=6432;
					out<=164;
				end
			end
			545: begin
				if(in == 0) begin
					state<=546;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=4444;
					out<=167;
				end
				if(in == 3) begin
					state<=2544;
					out<=168;
				end
				if(in == 4) begin
					state<=6433;
					out<=169;
				end
			end
			546: begin
				if(in == 0) begin
					state<=547;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=4445;
					out<=172;
				end
				if(in == 3) begin
					state<=2545;
					out<=173;
				end
				if(in == 4) begin
					state<=6434;
					out<=174;
				end
			end
			547: begin
				if(in == 0) begin
					state<=548;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=4446;
					out<=177;
				end
				if(in == 3) begin
					state<=2546;
					out<=178;
				end
				if(in == 4) begin
					state<=6435;
					out<=179;
				end
			end
			548: begin
				if(in == 0) begin
					state<=549;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=4447;
					out<=182;
				end
				if(in == 3) begin
					state<=2547;
					out<=183;
				end
				if(in == 4) begin
					state<=6436;
					out<=184;
				end
			end
			549: begin
				if(in == 0) begin
					state<=550;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=4448;
					out<=187;
				end
				if(in == 3) begin
					state<=2548;
					out<=188;
				end
				if(in == 4) begin
					state<=6437;
					out<=189;
				end
			end
			550: begin
				if(in == 0) begin
					state<=551;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=4449;
					out<=192;
				end
				if(in == 3) begin
					state<=2549;
					out<=193;
				end
				if(in == 4) begin
					state<=6438;
					out<=194;
				end
			end
			551: begin
				if(in == 0) begin
					state<=552;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=4450;
					out<=197;
				end
				if(in == 3) begin
					state<=2550;
					out<=198;
				end
				if(in == 4) begin
					state<=6439;
					out<=199;
				end
			end
			552: begin
				if(in == 0) begin
					state<=553;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=4451;
					out<=202;
				end
				if(in == 3) begin
					state<=2551;
					out<=203;
				end
				if(in == 4) begin
					state<=6440;
					out<=204;
				end
			end
			553: begin
				if(in == 0) begin
					state<=554;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=4452;
					out<=207;
				end
				if(in == 3) begin
					state<=2552;
					out<=208;
				end
				if(in == 4) begin
					state<=6441;
					out<=209;
				end
			end
			554: begin
				if(in == 0) begin
					state<=555;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=4453;
					out<=212;
				end
				if(in == 3) begin
					state<=2553;
					out<=213;
				end
				if(in == 4) begin
					state<=6442;
					out<=214;
				end
			end
			555: begin
				if(in == 0) begin
					state<=556;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=4454;
					out<=217;
				end
				if(in == 3) begin
					state<=2554;
					out<=218;
				end
				if(in == 4) begin
					state<=6443;
					out<=219;
				end
			end
			556: begin
				if(in == 0) begin
					state<=557;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=4455;
					out<=222;
				end
				if(in == 3) begin
					state<=2555;
					out<=223;
				end
				if(in == 4) begin
					state<=6444;
					out<=224;
				end
			end
			557: begin
				if(in == 0) begin
					state<=558;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=4456;
					out<=227;
				end
				if(in == 3) begin
					state<=2556;
					out<=228;
				end
				if(in == 4) begin
					state<=6445;
					out<=229;
				end
			end
			558: begin
				if(in == 0) begin
					state<=559;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=4457;
					out<=232;
				end
				if(in == 3) begin
					state<=2557;
					out<=233;
				end
				if(in == 4) begin
					state<=6446;
					out<=234;
				end
			end
			559: begin
				if(in == 0) begin
					state<=560;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=4458;
					out<=237;
				end
				if(in == 3) begin
					state<=2558;
					out<=238;
				end
				if(in == 4) begin
					state<=6447;
					out<=239;
				end
			end
			560: begin
				if(in == 0) begin
					state<=561;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=4459;
					out<=242;
				end
				if(in == 3) begin
					state<=2559;
					out<=243;
				end
				if(in == 4) begin
					state<=6448;
					out<=244;
				end
			end
			561: begin
				if(in == 0) begin
					state<=562;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=4460;
					out<=247;
				end
				if(in == 3) begin
					state<=2560;
					out<=248;
				end
				if(in == 4) begin
					state<=6449;
					out<=249;
				end
			end
			562: begin
				if(in == 0) begin
					state<=563;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=4461;
					out<=252;
				end
				if(in == 3) begin
					state<=2561;
					out<=253;
				end
				if(in == 4) begin
					state<=6450;
					out<=254;
				end
			end
			563: begin
				if(in == 0) begin
					state<=564;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=4462;
					out<=1;
				end
				if(in == 3) begin
					state<=2562;
					out<=2;
				end
				if(in == 4) begin
					state<=6451;
					out<=3;
				end
			end
			564: begin
				if(in == 0) begin
					state<=565;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=4463;
					out<=6;
				end
				if(in == 3) begin
					state<=2563;
					out<=7;
				end
				if(in == 4) begin
					state<=6452;
					out<=8;
				end
			end
			565: begin
				if(in == 0) begin
					state<=566;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=4464;
					out<=11;
				end
				if(in == 3) begin
					state<=2564;
					out<=12;
				end
				if(in == 4) begin
					state<=6453;
					out<=13;
				end
			end
			566: begin
				if(in == 0) begin
					state<=567;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=4465;
					out<=16;
				end
				if(in == 3) begin
					state<=2565;
					out<=17;
				end
				if(in == 4) begin
					state<=6454;
					out<=18;
				end
			end
			567: begin
				if(in == 0) begin
					state<=568;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=4466;
					out<=21;
				end
				if(in == 3) begin
					state<=2566;
					out<=22;
				end
				if(in == 4) begin
					state<=6455;
					out<=23;
				end
			end
			568: begin
				if(in == 0) begin
					state<=569;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=4467;
					out<=26;
				end
				if(in == 3) begin
					state<=2567;
					out<=27;
				end
				if(in == 4) begin
					state<=6456;
					out<=28;
				end
			end
			569: begin
				if(in == 0) begin
					state<=570;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=4468;
					out<=31;
				end
				if(in == 3) begin
					state<=2568;
					out<=32;
				end
				if(in == 4) begin
					state<=6457;
					out<=33;
				end
			end
			570: begin
				if(in == 0) begin
					state<=571;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=4469;
					out<=36;
				end
				if(in == 3) begin
					state<=2569;
					out<=37;
				end
				if(in == 4) begin
					state<=6458;
					out<=38;
				end
			end
			571: begin
				if(in == 0) begin
					state<=572;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=4470;
					out<=41;
				end
				if(in == 3) begin
					state<=2570;
					out<=42;
				end
				if(in == 4) begin
					state<=6459;
					out<=43;
				end
			end
			572: begin
				if(in == 0) begin
					state<=573;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=4471;
					out<=46;
				end
				if(in == 3) begin
					state<=2571;
					out<=47;
				end
				if(in == 4) begin
					state<=6460;
					out<=48;
				end
			end
			573: begin
				if(in == 0) begin
					state<=574;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=4472;
					out<=51;
				end
				if(in == 3) begin
					state<=2572;
					out<=52;
				end
				if(in == 4) begin
					state<=6461;
					out<=53;
				end
			end
			574: begin
				if(in == 0) begin
					state<=575;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=4473;
					out<=56;
				end
				if(in == 3) begin
					state<=2573;
					out<=57;
				end
				if(in == 4) begin
					state<=6462;
					out<=58;
				end
			end
			575: begin
				if(in == 0) begin
					state<=576;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=4474;
					out<=61;
				end
				if(in == 3) begin
					state<=2574;
					out<=62;
				end
				if(in == 4) begin
					state<=6463;
					out<=63;
				end
			end
			576: begin
				if(in == 0) begin
					state<=577;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=4475;
					out<=66;
				end
				if(in == 3) begin
					state<=2575;
					out<=67;
				end
				if(in == 4) begin
					state<=6464;
					out<=68;
				end
			end
			577: begin
				if(in == 0) begin
					state<=578;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=4476;
					out<=71;
				end
				if(in == 3) begin
					state<=2576;
					out<=72;
				end
				if(in == 4) begin
					state<=6465;
					out<=73;
				end
			end
			578: begin
				if(in == 0) begin
					state<=579;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=4477;
					out<=76;
				end
				if(in == 3) begin
					state<=2577;
					out<=77;
				end
				if(in == 4) begin
					state<=6466;
					out<=78;
				end
			end
			579: begin
				if(in == 0) begin
					state<=580;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=4478;
					out<=81;
				end
				if(in == 3) begin
					state<=2578;
					out<=82;
				end
				if(in == 4) begin
					state<=6467;
					out<=83;
				end
			end
			580: begin
				if(in == 0) begin
					state<=581;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=4479;
					out<=86;
				end
				if(in == 3) begin
					state<=2579;
					out<=87;
				end
				if(in == 4) begin
					state<=6468;
					out<=88;
				end
			end
			581: begin
				if(in == 0) begin
					state<=582;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=4480;
					out<=91;
				end
				if(in == 3) begin
					state<=2580;
					out<=92;
				end
				if(in == 4) begin
					state<=6469;
					out<=93;
				end
			end
			582: begin
				if(in == 0) begin
					state<=583;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=4481;
					out<=96;
				end
				if(in == 3) begin
					state<=2581;
					out<=97;
				end
				if(in == 4) begin
					state<=6470;
					out<=98;
				end
			end
			583: begin
				if(in == 0) begin
					state<=584;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=4482;
					out<=101;
				end
				if(in == 3) begin
					state<=2582;
					out<=102;
				end
				if(in == 4) begin
					state<=6471;
					out<=103;
				end
			end
			584: begin
				if(in == 0) begin
					state<=585;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=4483;
					out<=106;
				end
				if(in == 3) begin
					state<=2583;
					out<=107;
				end
				if(in == 4) begin
					state<=6472;
					out<=108;
				end
			end
			585: begin
				if(in == 0) begin
					state<=586;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=4484;
					out<=111;
				end
				if(in == 3) begin
					state<=2584;
					out<=112;
				end
				if(in == 4) begin
					state<=6473;
					out<=113;
				end
			end
			586: begin
				if(in == 0) begin
					state<=587;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=4485;
					out<=116;
				end
				if(in == 3) begin
					state<=2585;
					out<=117;
				end
				if(in == 4) begin
					state<=6474;
					out<=118;
				end
			end
			587: begin
				if(in == 0) begin
					state<=588;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=4486;
					out<=121;
				end
				if(in == 3) begin
					state<=2586;
					out<=122;
				end
				if(in == 4) begin
					state<=6475;
					out<=123;
				end
			end
			588: begin
				if(in == 0) begin
					state<=589;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=4487;
					out<=126;
				end
				if(in == 3) begin
					state<=2587;
					out<=127;
				end
				if(in == 4) begin
					state<=6476;
					out<=128;
				end
			end
			589: begin
				if(in == 0) begin
					state<=590;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=4488;
					out<=131;
				end
				if(in == 3) begin
					state<=2588;
					out<=132;
				end
				if(in == 4) begin
					state<=6477;
					out<=133;
				end
			end
			590: begin
				if(in == 0) begin
					state<=591;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=4489;
					out<=136;
				end
				if(in == 3) begin
					state<=2589;
					out<=137;
				end
				if(in == 4) begin
					state<=6478;
					out<=138;
				end
			end
			591: begin
				if(in == 0) begin
					state<=592;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=4490;
					out<=141;
				end
				if(in == 3) begin
					state<=2590;
					out<=142;
				end
				if(in == 4) begin
					state<=6479;
					out<=143;
				end
			end
			592: begin
				if(in == 0) begin
					state<=593;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=4491;
					out<=146;
				end
				if(in == 3) begin
					state<=2591;
					out<=147;
				end
				if(in == 4) begin
					state<=6480;
					out<=148;
				end
			end
			593: begin
				if(in == 0) begin
					state<=594;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=4492;
					out<=151;
				end
				if(in == 3) begin
					state<=2592;
					out<=152;
				end
				if(in == 4) begin
					state<=6481;
					out<=153;
				end
			end
			594: begin
				if(in == 0) begin
					state<=595;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=4493;
					out<=156;
				end
				if(in == 3) begin
					state<=2593;
					out<=157;
				end
				if(in == 4) begin
					state<=6482;
					out<=158;
				end
			end
			595: begin
				if(in == 0) begin
					state<=596;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=4494;
					out<=161;
				end
				if(in == 3) begin
					state<=2594;
					out<=162;
				end
				if(in == 4) begin
					state<=6483;
					out<=163;
				end
			end
			596: begin
				if(in == 0) begin
					state<=597;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=4495;
					out<=166;
				end
				if(in == 3) begin
					state<=2595;
					out<=167;
				end
				if(in == 4) begin
					state<=6484;
					out<=168;
				end
			end
			597: begin
				if(in == 0) begin
					state<=598;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=4496;
					out<=171;
				end
				if(in == 3) begin
					state<=2596;
					out<=172;
				end
				if(in == 4) begin
					state<=6485;
					out<=173;
				end
			end
			598: begin
				if(in == 0) begin
					state<=599;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=4497;
					out<=176;
				end
				if(in == 3) begin
					state<=2597;
					out<=177;
				end
				if(in == 4) begin
					state<=6486;
					out<=178;
				end
			end
			599: begin
				if(in == 0) begin
					state<=600;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=4498;
					out<=181;
				end
				if(in == 3) begin
					state<=2598;
					out<=182;
				end
				if(in == 4) begin
					state<=6487;
					out<=183;
				end
			end
			600: begin
				if(in == 0) begin
					state<=601;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=4499;
					out<=186;
				end
				if(in == 3) begin
					state<=2599;
					out<=187;
				end
				if(in == 4) begin
					state<=6488;
					out<=188;
				end
			end
			601: begin
				if(in == 0) begin
					state<=602;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=4500;
					out<=191;
				end
				if(in == 3) begin
					state<=2600;
					out<=192;
				end
				if(in == 4) begin
					state<=6489;
					out<=193;
				end
			end
			602: begin
				if(in == 0) begin
					state<=1546;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=5435;
					out<=196;
				end
				if(in == 3) begin
					state<=3478;
					out<=197;
				end
				if(in == 4) begin
					state<=7367;
					out<=198;
				end
			end
			603: begin
				if(in == 0) begin
					state<=604;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=4502;
					out<=201;
				end
				if(in == 3) begin
					state<=2602;
					out<=202;
				end
				if(in == 4) begin
					state<=6491;
					out<=203;
				end
			end
			604: begin
				if(in == 0) begin
					state<=605;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=4503;
					out<=206;
				end
				if(in == 3) begin
					state<=2603;
					out<=207;
				end
				if(in == 4) begin
					state<=6492;
					out<=208;
				end
			end
			605: begin
				if(in == 0) begin
					state<=606;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=4504;
					out<=211;
				end
				if(in == 3) begin
					state<=2604;
					out<=212;
				end
				if(in == 4) begin
					state<=6493;
					out<=213;
				end
			end
			606: begin
				if(in == 0) begin
					state<=607;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=4505;
					out<=216;
				end
				if(in == 3) begin
					state<=2605;
					out<=217;
				end
				if(in == 4) begin
					state<=6494;
					out<=218;
				end
			end
			607: begin
				if(in == 0) begin
					state<=608;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=4506;
					out<=221;
				end
				if(in == 3) begin
					state<=2606;
					out<=222;
				end
				if(in == 4) begin
					state<=6495;
					out<=223;
				end
			end
			608: begin
				if(in == 0) begin
					state<=609;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=4507;
					out<=226;
				end
				if(in == 3) begin
					state<=2607;
					out<=227;
				end
				if(in == 4) begin
					state<=6496;
					out<=228;
				end
			end
			609: begin
				if(in == 0) begin
					state<=610;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=4508;
					out<=231;
				end
				if(in == 3) begin
					state<=2608;
					out<=232;
				end
				if(in == 4) begin
					state<=6497;
					out<=233;
				end
			end
			610: begin
				if(in == 0) begin
					state<=611;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=4509;
					out<=236;
				end
				if(in == 3) begin
					state<=2609;
					out<=237;
				end
				if(in == 4) begin
					state<=6498;
					out<=238;
				end
			end
			611: begin
				if(in == 0) begin
					state<=612;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=4510;
					out<=241;
				end
				if(in == 3) begin
					state<=2610;
					out<=242;
				end
				if(in == 4) begin
					state<=6499;
					out<=243;
				end
			end
			612: begin
				if(in == 0) begin
					state<=613;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=4511;
					out<=246;
				end
				if(in == 3) begin
					state<=2611;
					out<=247;
				end
				if(in == 4) begin
					state<=6500;
					out<=248;
				end
			end
			613: begin
				if(in == 0) begin
					state<=614;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=4512;
					out<=251;
				end
				if(in == 3) begin
					state<=2612;
					out<=252;
				end
				if(in == 4) begin
					state<=6501;
					out<=253;
				end
			end
			614: begin
				if(in == 0) begin
					state<=615;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=4513;
					out<=0;
				end
				if(in == 3) begin
					state<=2613;
					out<=1;
				end
				if(in == 4) begin
					state<=6502;
					out<=2;
				end
			end
			615: begin
				if(in == 0) begin
					state<=616;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=4514;
					out<=5;
				end
				if(in == 3) begin
					state<=2614;
					out<=6;
				end
				if(in == 4) begin
					state<=6503;
					out<=7;
				end
			end
			616: begin
				if(in == 0) begin
					state<=617;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=4515;
					out<=10;
				end
				if(in == 3) begin
					state<=2615;
					out<=11;
				end
				if(in == 4) begin
					state<=6504;
					out<=12;
				end
			end
			617: begin
				if(in == 0) begin
					state<=618;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=4516;
					out<=15;
				end
				if(in == 3) begin
					state<=2616;
					out<=16;
				end
				if(in == 4) begin
					state<=6505;
					out<=17;
				end
			end
			618: begin
				if(in == 0) begin
					state<=619;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=4517;
					out<=20;
				end
				if(in == 3) begin
					state<=2617;
					out<=21;
				end
				if(in == 4) begin
					state<=6506;
					out<=22;
				end
			end
			619: begin
				if(in == 0) begin
					state<=620;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=4518;
					out<=25;
				end
				if(in == 3) begin
					state<=2618;
					out<=26;
				end
				if(in == 4) begin
					state<=6507;
					out<=27;
				end
			end
			620: begin
				if(in == 0) begin
					state<=621;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=4519;
					out<=30;
				end
				if(in == 3) begin
					state<=2619;
					out<=31;
				end
				if(in == 4) begin
					state<=6508;
					out<=32;
				end
			end
			621: begin
				if(in == 0) begin
					state<=622;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=4520;
					out<=35;
				end
				if(in == 3) begin
					state<=2620;
					out<=36;
				end
				if(in == 4) begin
					state<=6509;
					out<=37;
				end
			end
			622: begin
				if(in == 0) begin
					state<=623;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=4521;
					out<=40;
				end
				if(in == 3) begin
					state<=2621;
					out<=41;
				end
				if(in == 4) begin
					state<=6510;
					out<=42;
				end
			end
			623: begin
				if(in == 0) begin
					state<=624;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=4522;
					out<=45;
				end
				if(in == 3) begin
					state<=2622;
					out<=46;
				end
				if(in == 4) begin
					state<=6511;
					out<=47;
				end
			end
			624: begin
				if(in == 0) begin
					state<=625;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=4523;
					out<=50;
				end
				if(in == 3) begin
					state<=2623;
					out<=51;
				end
				if(in == 4) begin
					state<=6512;
					out<=52;
				end
			end
			625: begin
				if(in == 0) begin
					state<=626;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=4524;
					out<=55;
				end
				if(in == 3) begin
					state<=2624;
					out<=56;
				end
				if(in == 4) begin
					state<=6513;
					out<=57;
				end
			end
			626: begin
				if(in == 0) begin
					state<=627;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=4525;
					out<=60;
				end
				if(in == 3) begin
					state<=2625;
					out<=61;
				end
				if(in == 4) begin
					state<=6514;
					out<=62;
				end
			end
			627: begin
				if(in == 0) begin
					state<=628;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=4526;
					out<=65;
				end
				if(in == 3) begin
					state<=2626;
					out<=66;
				end
				if(in == 4) begin
					state<=6515;
					out<=67;
				end
			end
			628: begin
				if(in == 0) begin
					state<=629;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=4527;
					out<=70;
				end
				if(in == 3) begin
					state<=2627;
					out<=71;
				end
				if(in == 4) begin
					state<=6516;
					out<=72;
				end
			end
			629: begin
				if(in == 0) begin
					state<=630;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=4528;
					out<=75;
				end
				if(in == 3) begin
					state<=2628;
					out<=76;
				end
				if(in == 4) begin
					state<=6517;
					out<=77;
				end
			end
			630: begin
				if(in == 0) begin
					state<=631;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=4529;
					out<=80;
				end
				if(in == 3) begin
					state<=2629;
					out<=81;
				end
				if(in == 4) begin
					state<=6518;
					out<=82;
				end
			end
			631: begin
				if(in == 0) begin
					state<=632;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=4530;
					out<=85;
				end
				if(in == 3) begin
					state<=2630;
					out<=86;
				end
				if(in == 4) begin
					state<=6519;
					out<=87;
				end
			end
			632: begin
				if(in == 0) begin
					state<=633;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=4531;
					out<=90;
				end
				if(in == 3) begin
					state<=2631;
					out<=91;
				end
				if(in == 4) begin
					state<=6520;
					out<=92;
				end
			end
			633: begin
				if(in == 0) begin
					state<=634;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=4532;
					out<=95;
				end
				if(in == 3) begin
					state<=2632;
					out<=96;
				end
				if(in == 4) begin
					state<=6521;
					out<=97;
				end
			end
			634: begin
				if(in == 0) begin
					state<=635;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=4533;
					out<=100;
				end
				if(in == 3) begin
					state<=2633;
					out<=101;
				end
				if(in == 4) begin
					state<=6522;
					out<=102;
				end
			end
			635: begin
				if(in == 0) begin
					state<=636;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=4534;
					out<=105;
				end
				if(in == 3) begin
					state<=2634;
					out<=106;
				end
				if(in == 4) begin
					state<=6523;
					out<=107;
				end
			end
			636: begin
				if(in == 0) begin
					state<=637;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=4535;
					out<=110;
				end
				if(in == 3) begin
					state<=2635;
					out<=111;
				end
				if(in == 4) begin
					state<=6524;
					out<=112;
				end
			end
			637: begin
				if(in == 0) begin
					state<=638;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=4536;
					out<=115;
				end
				if(in == 3) begin
					state<=2636;
					out<=116;
				end
				if(in == 4) begin
					state<=6525;
					out<=117;
				end
			end
			638: begin
				if(in == 0) begin
					state<=639;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=4537;
					out<=120;
				end
				if(in == 3) begin
					state<=2637;
					out<=121;
				end
				if(in == 4) begin
					state<=6526;
					out<=122;
				end
			end
			639: begin
				if(in == 0) begin
					state<=640;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=4538;
					out<=125;
				end
				if(in == 3) begin
					state<=2638;
					out<=126;
				end
				if(in == 4) begin
					state<=6527;
					out<=127;
				end
			end
			640: begin
				if(in == 0) begin
					state<=641;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=4539;
					out<=130;
				end
				if(in == 3) begin
					state<=2639;
					out<=131;
				end
				if(in == 4) begin
					state<=6528;
					out<=132;
				end
			end
			641: begin
				if(in == 0) begin
					state<=642;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=4540;
					out<=135;
				end
				if(in == 3) begin
					state<=2640;
					out<=136;
				end
				if(in == 4) begin
					state<=6529;
					out<=137;
				end
			end
			642: begin
				if(in == 0) begin
					state<=643;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=4541;
					out<=140;
				end
				if(in == 3) begin
					state<=2641;
					out<=141;
				end
				if(in == 4) begin
					state<=6530;
					out<=142;
				end
			end
			643: begin
				if(in == 0) begin
					state<=644;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=4542;
					out<=145;
				end
				if(in == 3) begin
					state<=2642;
					out<=146;
				end
				if(in == 4) begin
					state<=6531;
					out<=147;
				end
			end
			644: begin
				if(in == 0) begin
					state<=645;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=4543;
					out<=150;
				end
				if(in == 3) begin
					state<=2643;
					out<=151;
				end
				if(in == 4) begin
					state<=6532;
					out<=152;
				end
			end
			645: begin
				if(in == 0) begin
					state<=646;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=4544;
					out<=155;
				end
				if(in == 3) begin
					state<=2644;
					out<=156;
				end
				if(in == 4) begin
					state<=6533;
					out<=157;
				end
			end
			646: begin
				if(in == 0) begin
					state<=647;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=4545;
					out<=160;
				end
				if(in == 3) begin
					state<=2645;
					out<=161;
				end
				if(in == 4) begin
					state<=6534;
					out<=162;
				end
			end
			647: begin
				if(in == 0) begin
					state<=648;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=4546;
					out<=165;
				end
				if(in == 3) begin
					state<=2646;
					out<=166;
				end
				if(in == 4) begin
					state<=6535;
					out<=167;
				end
			end
			648: begin
				if(in == 0) begin
					state<=649;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=4547;
					out<=170;
				end
				if(in == 3) begin
					state<=2647;
					out<=171;
				end
				if(in == 4) begin
					state<=6536;
					out<=172;
				end
			end
			649: begin
				if(in == 0) begin
					state<=650;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=4548;
					out<=175;
				end
				if(in == 3) begin
					state<=2648;
					out<=176;
				end
				if(in == 4) begin
					state<=6537;
					out<=177;
				end
			end
			650: begin
				if(in == 0) begin
					state<=651;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=4549;
					out<=180;
				end
				if(in == 3) begin
					state<=2649;
					out<=181;
				end
				if(in == 4) begin
					state<=6538;
					out<=182;
				end
			end
			651: begin
				if(in == 0) begin
					state<=652;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=4550;
					out<=185;
				end
				if(in == 3) begin
					state<=2650;
					out<=186;
				end
				if(in == 4) begin
					state<=6539;
					out<=187;
				end
			end
			652: begin
				if(in == 0) begin
					state<=653;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=4551;
					out<=190;
				end
				if(in == 3) begin
					state<=2651;
					out<=191;
				end
				if(in == 4) begin
					state<=6540;
					out<=192;
				end
			end
			653: begin
				if(in == 0) begin
					state<=654;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=4552;
					out<=195;
				end
				if(in == 3) begin
					state<=2652;
					out<=196;
				end
				if(in == 4) begin
					state<=6541;
					out<=197;
				end
			end
			654: begin
				if(in == 0) begin
					state<=655;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=4553;
					out<=200;
				end
				if(in == 3) begin
					state<=2653;
					out<=201;
				end
				if(in == 4) begin
					state<=6542;
					out<=202;
				end
			end
			655: begin
				if(in == 0) begin
					state<=656;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=4554;
					out<=205;
				end
				if(in == 3) begin
					state<=2654;
					out<=206;
				end
				if(in == 4) begin
					state<=6543;
					out<=207;
				end
			end
			656: begin
				if(in == 0) begin
					state<=657;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=4555;
					out<=210;
				end
				if(in == 3) begin
					state<=2655;
					out<=211;
				end
				if(in == 4) begin
					state<=6544;
					out<=212;
				end
			end
			657: begin
				if(in == 0) begin
					state<=658;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=4556;
					out<=215;
				end
				if(in == 3) begin
					state<=2656;
					out<=216;
				end
				if(in == 4) begin
					state<=6545;
					out<=217;
				end
			end
			658: begin
				if(in == 0) begin
					state<=659;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=4557;
					out<=220;
				end
				if(in == 3) begin
					state<=2657;
					out<=221;
				end
				if(in == 4) begin
					state<=6546;
					out<=222;
				end
			end
			659: begin
				if(in == 0) begin
					state<=660;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=4558;
					out<=225;
				end
				if(in == 3) begin
					state<=2658;
					out<=226;
				end
				if(in == 4) begin
					state<=6547;
					out<=227;
				end
			end
			660: begin
				if(in == 0) begin
					state<=661;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=4559;
					out<=230;
				end
				if(in == 3) begin
					state<=2659;
					out<=231;
				end
				if(in == 4) begin
					state<=6548;
					out<=232;
				end
			end
			661: begin
				if(in == 0) begin
					state<=662;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=4560;
					out<=235;
				end
				if(in == 3) begin
					state<=2660;
					out<=236;
				end
				if(in == 4) begin
					state<=6549;
					out<=237;
				end
			end
			662: begin
				if(in == 0) begin
					state<=663;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=4561;
					out<=240;
				end
				if(in == 3) begin
					state<=2661;
					out<=241;
				end
				if(in == 4) begin
					state<=6550;
					out<=242;
				end
			end
			663: begin
				if(in == 0) begin
					state<=664;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=4562;
					out<=245;
				end
				if(in == 3) begin
					state<=2662;
					out<=246;
				end
				if(in == 4) begin
					state<=6551;
					out<=247;
				end
			end
			664: begin
				if(in == 0) begin
					state<=665;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=4563;
					out<=250;
				end
				if(in == 3) begin
					state<=2663;
					out<=251;
				end
				if(in == 4) begin
					state<=6552;
					out<=252;
				end
			end
			665: begin
				if(in == 0) begin
					state<=666;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=4564;
					out<=255;
				end
				if(in == 3) begin
					state<=2664;
					out<=0;
				end
				if(in == 4) begin
					state<=6553;
					out<=1;
				end
			end
			666: begin
				if(in == 0) begin
					state<=667;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=4565;
					out<=4;
				end
				if(in == 3) begin
					state<=2665;
					out<=5;
				end
				if(in == 4) begin
					state<=6554;
					out<=6;
				end
			end
			667: begin
				if(in == 0) begin
					state<=668;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=4566;
					out<=9;
				end
				if(in == 3) begin
					state<=2666;
					out<=10;
				end
				if(in == 4) begin
					state<=6555;
					out<=11;
				end
			end
			668: begin
				if(in == 0) begin
					state<=669;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=4567;
					out<=14;
				end
				if(in == 3) begin
					state<=2667;
					out<=15;
				end
				if(in == 4) begin
					state<=6556;
					out<=16;
				end
			end
			669: begin
				if(in == 0) begin
					state<=670;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=4568;
					out<=19;
				end
				if(in == 3) begin
					state<=2668;
					out<=20;
				end
				if(in == 4) begin
					state<=6557;
					out<=21;
				end
			end
			670: begin
				if(in == 0) begin
					state<=671;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=4569;
					out<=24;
				end
				if(in == 3) begin
					state<=2669;
					out<=25;
				end
				if(in == 4) begin
					state<=6558;
					out<=26;
				end
			end
			671: begin
				if(in == 0) begin
					state<=1577;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=5466;
					out<=29;
				end
				if(in == 3) begin
					state<=3230;
					out<=30;
				end
				if(in == 4) begin
					state<=7119;
					out<=31;
				end
			end
			672: begin
				if(in == 0) begin
					state<=673;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=4571;
					out<=34;
				end
				if(in == 3) begin
					state<=2671;
					out<=35;
				end
				if(in == 4) begin
					state<=6560;
					out<=36;
				end
			end
			673: begin
				if(in == 0) begin
					state<=674;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=4572;
					out<=39;
				end
				if(in == 3) begin
					state<=2672;
					out<=40;
				end
				if(in == 4) begin
					state<=6561;
					out<=41;
				end
			end
			674: begin
				if(in == 0) begin
					state<=675;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=4573;
					out<=44;
				end
				if(in == 3) begin
					state<=2673;
					out<=45;
				end
				if(in == 4) begin
					state<=6562;
					out<=46;
				end
			end
			675: begin
				if(in == 0) begin
					state<=676;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=4574;
					out<=49;
				end
				if(in == 3) begin
					state<=2674;
					out<=50;
				end
				if(in == 4) begin
					state<=6563;
					out<=51;
				end
			end
			676: begin
				if(in == 0) begin
					state<=677;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=4575;
					out<=54;
				end
				if(in == 3) begin
					state<=2675;
					out<=55;
				end
				if(in == 4) begin
					state<=6564;
					out<=56;
				end
			end
			677: begin
				if(in == 0) begin
					state<=678;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=4576;
					out<=59;
				end
				if(in == 3) begin
					state<=2676;
					out<=60;
				end
				if(in == 4) begin
					state<=6565;
					out<=61;
				end
			end
			678: begin
				if(in == 0) begin
					state<=679;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=4577;
					out<=64;
				end
				if(in == 3) begin
					state<=2677;
					out<=65;
				end
				if(in == 4) begin
					state<=6566;
					out<=66;
				end
			end
			679: begin
				if(in == 0) begin
					state<=680;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=4578;
					out<=69;
				end
				if(in == 3) begin
					state<=2678;
					out<=70;
				end
				if(in == 4) begin
					state<=6567;
					out<=71;
				end
			end
			680: begin
				if(in == 0) begin
					state<=681;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=4579;
					out<=74;
				end
				if(in == 3) begin
					state<=2679;
					out<=75;
				end
				if(in == 4) begin
					state<=6568;
					out<=76;
				end
			end
			681: begin
				if(in == 0) begin
					state<=682;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=4580;
					out<=79;
				end
				if(in == 3) begin
					state<=2680;
					out<=80;
				end
				if(in == 4) begin
					state<=6569;
					out<=81;
				end
			end
			682: begin
				if(in == 0) begin
					state<=683;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=4581;
					out<=84;
				end
				if(in == 3) begin
					state<=2681;
					out<=85;
				end
				if(in == 4) begin
					state<=6570;
					out<=86;
				end
			end
			683: begin
				if(in == 0) begin
					state<=684;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=4582;
					out<=89;
				end
				if(in == 3) begin
					state<=2682;
					out<=90;
				end
				if(in == 4) begin
					state<=6571;
					out<=91;
				end
			end
			684: begin
				if(in == 0) begin
					state<=685;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=4583;
					out<=94;
				end
				if(in == 3) begin
					state<=2683;
					out<=95;
				end
				if(in == 4) begin
					state<=6572;
					out<=96;
				end
			end
			685: begin
				if(in == 0) begin
					state<=686;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=4584;
					out<=99;
				end
				if(in == 3) begin
					state<=2684;
					out<=100;
				end
				if(in == 4) begin
					state<=6573;
					out<=101;
				end
			end
			686: begin
				if(in == 0) begin
					state<=687;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=4585;
					out<=104;
				end
				if(in == 3) begin
					state<=2685;
					out<=105;
				end
				if(in == 4) begin
					state<=6574;
					out<=106;
				end
			end
			687: begin
				if(in == 0) begin
					state<=688;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=4586;
					out<=109;
				end
				if(in == 3) begin
					state<=2686;
					out<=110;
				end
				if(in == 4) begin
					state<=6575;
					out<=111;
				end
			end
			688: begin
				if(in == 0) begin
					state<=689;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=4587;
					out<=114;
				end
				if(in == 3) begin
					state<=2687;
					out<=115;
				end
				if(in == 4) begin
					state<=6576;
					out<=116;
				end
			end
			689: begin
				if(in == 0) begin
					state<=690;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=4588;
					out<=119;
				end
				if(in == 3) begin
					state<=2688;
					out<=120;
				end
				if(in == 4) begin
					state<=6577;
					out<=121;
				end
			end
			690: begin
				if(in == 0) begin
					state<=1;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=3899;
					out<=124;
				end
				if(in == 3) begin
					state<=1999;
					out<=125;
				end
				if(in == 4) begin
					state<=5888;
					out<=126;
				end
			end
			691: begin
				if(in == 0) begin
					state<=692;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=4590;
					out<=129;
				end
				if(in == 3) begin
					state<=2690;
					out<=130;
				end
				if(in == 4) begin
					state<=6579;
					out<=131;
				end
			end
			692: begin
				if(in == 0) begin
					state<=693;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=4591;
					out<=134;
				end
				if(in == 3) begin
					state<=2691;
					out<=135;
				end
				if(in == 4) begin
					state<=6580;
					out<=136;
				end
			end
			693: begin
				if(in == 0) begin
					state<=694;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=4592;
					out<=139;
				end
				if(in == 3) begin
					state<=2692;
					out<=140;
				end
				if(in == 4) begin
					state<=6581;
					out<=141;
				end
			end
			694: begin
				if(in == 0) begin
					state<=695;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=4593;
					out<=144;
				end
				if(in == 3) begin
					state<=2693;
					out<=145;
				end
				if(in == 4) begin
					state<=6582;
					out<=146;
				end
			end
			695: begin
				if(in == 0) begin
					state<=696;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=4594;
					out<=149;
				end
				if(in == 3) begin
					state<=2694;
					out<=150;
				end
				if(in == 4) begin
					state<=6583;
					out<=151;
				end
			end
			696: begin
				if(in == 0) begin
					state<=697;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=4595;
					out<=154;
				end
				if(in == 3) begin
					state<=2695;
					out<=155;
				end
				if(in == 4) begin
					state<=6584;
					out<=156;
				end
			end
			697: begin
				if(in == 0) begin
					state<=698;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=4596;
					out<=159;
				end
				if(in == 3) begin
					state<=2696;
					out<=160;
				end
				if(in == 4) begin
					state<=6585;
					out<=161;
				end
			end
			698: begin
				if(in == 0) begin
					state<=699;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=4597;
					out<=164;
				end
				if(in == 3) begin
					state<=2697;
					out<=165;
				end
				if(in == 4) begin
					state<=6586;
					out<=166;
				end
			end
			699: begin
				if(in == 0) begin
					state<=700;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=4598;
					out<=169;
				end
				if(in == 3) begin
					state<=2698;
					out<=170;
				end
				if(in == 4) begin
					state<=6587;
					out<=171;
				end
			end
			700: begin
				if(in == 0) begin
					state<=701;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=4599;
					out<=174;
				end
				if(in == 3) begin
					state<=2699;
					out<=175;
				end
				if(in == 4) begin
					state<=6588;
					out<=176;
				end
			end
			701: begin
				if(in == 0) begin
					state<=702;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=4600;
					out<=179;
				end
				if(in == 3) begin
					state<=2700;
					out<=180;
				end
				if(in == 4) begin
					state<=6589;
					out<=181;
				end
			end
			702: begin
				if(in == 0) begin
					state<=703;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=4601;
					out<=184;
				end
				if(in == 3) begin
					state<=2701;
					out<=185;
				end
				if(in == 4) begin
					state<=6590;
					out<=186;
				end
			end
			703: begin
				if(in == 0) begin
					state<=704;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=4602;
					out<=189;
				end
				if(in == 3) begin
					state<=2702;
					out<=190;
				end
				if(in == 4) begin
					state<=6591;
					out<=191;
				end
			end
			704: begin
				if(in == 0) begin
					state<=705;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=4603;
					out<=194;
				end
				if(in == 3) begin
					state<=2703;
					out<=195;
				end
				if(in == 4) begin
					state<=6592;
					out<=196;
				end
			end
			705: begin
				if(in == 0) begin
					state<=706;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=4604;
					out<=199;
				end
				if(in == 3) begin
					state<=2704;
					out<=200;
				end
				if(in == 4) begin
					state<=6593;
					out<=201;
				end
			end
			706: begin
				if(in == 0) begin
					state<=707;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=4605;
					out<=204;
				end
				if(in == 3) begin
					state<=2705;
					out<=205;
				end
				if(in == 4) begin
					state<=6594;
					out<=206;
				end
			end
			707: begin
				if(in == 0) begin
					state<=708;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=4606;
					out<=209;
				end
				if(in == 3) begin
					state<=2706;
					out<=210;
				end
				if(in == 4) begin
					state<=6595;
					out<=211;
				end
			end
			708: begin
				if(in == 0) begin
					state<=709;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=4607;
					out<=214;
				end
				if(in == 3) begin
					state<=2707;
					out<=215;
				end
				if(in == 4) begin
					state<=6596;
					out<=216;
				end
			end
			709: begin
				if(in == 0) begin
					state<=710;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=4608;
					out<=219;
				end
				if(in == 3) begin
					state<=2708;
					out<=220;
				end
				if(in == 4) begin
					state<=6597;
					out<=221;
				end
			end
			710: begin
				if(in == 0) begin
					state<=711;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=4609;
					out<=224;
				end
				if(in == 3) begin
					state<=2709;
					out<=225;
				end
				if(in == 4) begin
					state<=6598;
					out<=226;
				end
			end
			711: begin
				if(in == 0) begin
					state<=712;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=4610;
					out<=229;
				end
				if(in == 3) begin
					state<=2710;
					out<=230;
				end
				if(in == 4) begin
					state<=6599;
					out<=231;
				end
			end
			712: begin
				if(in == 0) begin
					state<=713;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=4611;
					out<=234;
				end
				if(in == 3) begin
					state<=2711;
					out<=235;
				end
				if(in == 4) begin
					state<=6600;
					out<=236;
				end
			end
			713: begin
				if(in == 0) begin
					state<=714;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=4612;
					out<=239;
				end
				if(in == 3) begin
					state<=2712;
					out<=240;
				end
				if(in == 4) begin
					state<=6601;
					out<=241;
				end
			end
			714: begin
				if(in == 0) begin
					state<=715;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=4613;
					out<=244;
				end
				if(in == 3) begin
					state<=2713;
					out<=245;
				end
				if(in == 4) begin
					state<=6602;
					out<=246;
				end
			end
			715: begin
				if(in == 0) begin
					state<=716;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=4614;
					out<=249;
				end
				if(in == 3) begin
					state<=2714;
					out<=250;
				end
				if(in == 4) begin
					state<=6603;
					out<=251;
				end
			end
			716: begin
				if(in == 0) begin
					state<=717;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=4615;
					out<=254;
				end
				if(in == 3) begin
					state<=2715;
					out<=255;
				end
				if(in == 4) begin
					state<=6604;
					out<=0;
				end
			end
			717: begin
				if(in == 0) begin
					state<=718;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=4616;
					out<=3;
				end
				if(in == 3) begin
					state<=2716;
					out<=4;
				end
				if(in == 4) begin
					state<=6605;
					out<=5;
				end
			end
			718: begin
				if(in == 0) begin
					state<=719;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=4617;
					out<=8;
				end
				if(in == 3) begin
					state<=2717;
					out<=9;
				end
				if(in == 4) begin
					state<=6606;
					out<=10;
				end
			end
			719: begin
				if(in == 0) begin
					state<=720;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=4618;
					out<=13;
				end
				if(in == 3) begin
					state<=2718;
					out<=14;
				end
				if(in == 4) begin
					state<=6607;
					out<=15;
				end
			end
			720: begin
				if(in == 0) begin
					state<=721;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=4619;
					out<=18;
				end
				if(in == 3) begin
					state<=2719;
					out<=19;
				end
				if(in == 4) begin
					state<=6608;
					out<=20;
				end
			end
			721: begin
				if(in == 0) begin
					state<=722;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=4620;
					out<=23;
				end
				if(in == 3) begin
					state<=2720;
					out<=24;
				end
				if(in == 4) begin
					state<=6609;
					out<=25;
				end
			end
			722: begin
				if(in == 0) begin
					state<=723;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=4621;
					out<=28;
				end
				if(in == 3) begin
					state<=2721;
					out<=29;
				end
				if(in == 4) begin
					state<=6610;
					out<=30;
				end
			end
			723: begin
				if(in == 0) begin
					state<=724;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=4622;
					out<=33;
				end
				if(in == 3) begin
					state<=2722;
					out<=34;
				end
				if(in == 4) begin
					state<=6611;
					out<=35;
				end
			end
			724: begin
				if(in == 0) begin
					state<=725;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=4623;
					out<=38;
				end
				if(in == 3) begin
					state<=2723;
					out<=39;
				end
				if(in == 4) begin
					state<=6612;
					out<=40;
				end
			end
			725: begin
				if(in == 0) begin
					state<=726;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=4624;
					out<=43;
				end
				if(in == 3) begin
					state<=2724;
					out<=44;
				end
				if(in == 4) begin
					state<=6613;
					out<=45;
				end
			end
			726: begin
				if(in == 0) begin
					state<=727;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=4625;
					out<=48;
				end
				if(in == 3) begin
					state<=2725;
					out<=49;
				end
				if(in == 4) begin
					state<=6614;
					out<=50;
				end
			end
			727: begin
				if(in == 0) begin
					state<=728;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=4626;
					out<=53;
				end
				if(in == 3) begin
					state<=2726;
					out<=54;
				end
				if(in == 4) begin
					state<=6615;
					out<=55;
				end
			end
			728: begin
				if(in == 0) begin
					state<=729;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=4627;
					out<=58;
				end
				if(in == 3) begin
					state<=2727;
					out<=59;
				end
				if(in == 4) begin
					state<=6616;
					out<=60;
				end
			end
			729: begin
				if(in == 0) begin
					state<=730;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=4628;
					out<=63;
				end
				if(in == 3) begin
					state<=2728;
					out<=64;
				end
				if(in == 4) begin
					state<=6617;
					out<=65;
				end
			end
			730: begin
				if(in == 0) begin
					state<=731;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=4629;
					out<=68;
				end
				if(in == 3) begin
					state<=2729;
					out<=69;
				end
				if(in == 4) begin
					state<=6618;
					out<=70;
				end
			end
			731: begin
				if(in == 0) begin
					state<=732;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=4630;
					out<=73;
				end
				if(in == 3) begin
					state<=2730;
					out<=74;
				end
				if(in == 4) begin
					state<=6619;
					out<=75;
				end
			end
			732: begin
				if(in == 0) begin
					state<=733;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=4631;
					out<=78;
				end
				if(in == 3) begin
					state<=2731;
					out<=79;
				end
				if(in == 4) begin
					state<=6620;
					out<=80;
				end
			end
			733: begin
				if(in == 0) begin
					state<=734;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=4632;
					out<=83;
				end
				if(in == 3) begin
					state<=2732;
					out<=84;
				end
				if(in == 4) begin
					state<=6621;
					out<=85;
				end
			end
			734: begin
				if(in == 0) begin
					state<=735;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=4633;
					out<=88;
				end
				if(in == 3) begin
					state<=2733;
					out<=89;
				end
				if(in == 4) begin
					state<=6622;
					out<=90;
				end
			end
			735: begin
				if(in == 0) begin
					state<=736;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=4634;
					out<=93;
				end
				if(in == 3) begin
					state<=2734;
					out<=94;
				end
				if(in == 4) begin
					state<=6623;
					out<=95;
				end
			end
			736: begin
				if(in == 0) begin
					state<=737;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=4635;
					out<=98;
				end
				if(in == 3) begin
					state<=2735;
					out<=99;
				end
				if(in == 4) begin
					state<=6624;
					out<=100;
				end
			end
			737: begin
				if(in == 0) begin
					state<=738;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=4636;
					out<=103;
				end
				if(in == 3) begin
					state<=2736;
					out<=104;
				end
				if(in == 4) begin
					state<=6625;
					out<=105;
				end
			end
			738: begin
				if(in == 0) begin
					state<=739;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=4637;
					out<=108;
				end
				if(in == 3) begin
					state<=2737;
					out<=109;
				end
				if(in == 4) begin
					state<=6626;
					out<=110;
				end
			end
			739: begin
				if(in == 0) begin
					state<=740;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=4638;
					out<=113;
				end
				if(in == 3) begin
					state<=2738;
					out<=114;
				end
				if(in == 4) begin
					state<=6627;
					out<=115;
				end
			end
			740: begin
				if(in == 0) begin
					state<=741;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=4639;
					out<=118;
				end
				if(in == 3) begin
					state<=2739;
					out<=119;
				end
				if(in == 4) begin
					state<=6628;
					out<=120;
				end
			end
			741: begin
				if(in == 0) begin
					state<=742;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=4640;
					out<=123;
				end
				if(in == 3) begin
					state<=2740;
					out<=124;
				end
				if(in == 4) begin
					state<=6629;
					out<=125;
				end
			end
			742: begin
				if(in == 0) begin
					state<=743;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=4641;
					out<=128;
				end
				if(in == 3) begin
					state<=2741;
					out<=129;
				end
				if(in == 4) begin
					state<=6630;
					out<=130;
				end
			end
			743: begin
				if(in == 0) begin
					state<=744;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=4642;
					out<=133;
				end
				if(in == 3) begin
					state<=2742;
					out<=134;
				end
				if(in == 4) begin
					state<=6631;
					out<=135;
				end
			end
			744: begin
				if(in == 0) begin
					state<=745;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=4643;
					out<=138;
				end
				if(in == 3) begin
					state<=2743;
					out<=139;
				end
				if(in == 4) begin
					state<=6632;
					out<=140;
				end
			end
			745: begin
				if(in == 0) begin
					state<=746;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=4644;
					out<=143;
				end
				if(in == 3) begin
					state<=2744;
					out<=144;
				end
				if(in == 4) begin
					state<=6633;
					out<=145;
				end
			end
			746: begin
				if(in == 0) begin
					state<=747;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=4645;
					out<=148;
				end
				if(in == 3) begin
					state<=2745;
					out<=149;
				end
				if(in == 4) begin
					state<=6634;
					out<=150;
				end
			end
			747: begin
				if(in == 0) begin
					state<=748;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=4646;
					out<=153;
				end
				if(in == 3) begin
					state<=2746;
					out<=154;
				end
				if(in == 4) begin
					state<=6635;
					out<=155;
				end
			end
			748: begin
				if(in == 0) begin
					state<=749;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=4647;
					out<=158;
				end
				if(in == 3) begin
					state<=2747;
					out<=159;
				end
				if(in == 4) begin
					state<=6636;
					out<=160;
				end
			end
			749: begin
				if(in == 0) begin
					state<=750;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=4648;
					out<=163;
				end
				if(in == 3) begin
					state<=2748;
					out<=164;
				end
				if(in == 4) begin
					state<=6637;
					out<=165;
				end
			end
			750: begin
				if(in == 0) begin
					state<=751;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=4649;
					out<=168;
				end
				if(in == 3) begin
					state<=2749;
					out<=169;
				end
				if(in == 4) begin
					state<=6638;
					out<=170;
				end
			end
			751: begin
				if(in == 0) begin
					state<=752;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=4650;
					out<=173;
				end
				if(in == 3) begin
					state<=2750;
					out<=174;
				end
				if(in == 4) begin
					state<=6639;
					out<=175;
				end
			end
			752: begin
				if(in == 0) begin
					state<=753;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=4651;
					out<=178;
				end
				if(in == 3) begin
					state<=2751;
					out<=179;
				end
				if(in == 4) begin
					state<=6640;
					out<=180;
				end
			end
			753: begin
				if(in == 0) begin
					state<=754;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=4652;
					out<=183;
				end
				if(in == 3) begin
					state<=2752;
					out<=184;
				end
				if(in == 4) begin
					state<=6641;
					out<=185;
				end
			end
			754: begin
				if(in == 0) begin
					state<=755;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=4653;
					out<=188;
				end
				if(in == 3) begin
					state<=2753;
					out<=189;
				end
				if(in == 4) begin
					state<=6642;
					out<=190;
				end
			end
			755: begin
				if(in == 0) begin
					state<=756;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=4654;
					out<=193;
				end
				if(in == 3) begin
					state<=2754;
					out<=194;
				end
				if(in == 4) begin
					state<=6643;
					out<=195;
				end
			end
			756: begin
				if(in == 0) begin
					state<=757;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=4655;
					out<=198;
				end
				if(in == 3) begin
					state<=2755;
					out<=199;
				end
				if(in == 4) begin
					state<=6644;
					out<=200;
				end
			end
			757: begin
				if(in == 0) begin
					state<=758;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=4656;
					out<=203;
				end
				if(in == 3) begin
					state<=2756;
					out<=204;
				end
				if(in == 4) begin
					state<=6645;
					out<=205;
				end
			end
			758: begin
				if(in == 0) begin
					state<=759;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=4657;
					out<=208;
				end
				if(in == 3) begin
					state<=2757;
					out<=209;
				end
				if(in == 4) begin
					state<=6646;
					out<=210;
				end
			end
			759: begin
				if(in == 0) begin
					state<=760;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=4658;
					out<=213;
				end
				if(in == 3) begin
					state<=2758;
					out<=214;
				end
				if(in == 4) begin
					state<=6647;
					out<=215;
				end
			end
			760: begin
				if(in == 0) begin
					state<=761;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=4659;
					out<=218;
				end
				if(in == 3) begin
					state<=2759;
					out<=219;
				end
				if(in == 4) begin
					state<=6648;
					out<=220;
				end
			end
			761: begin
				if(in == 0) begin
					state<=762;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=4660;
					out<=223;
				end
				if(in == 3) begin
					state<=2760;
					out<=224;
				end
				if(in == 4) begin
					state<=6649;
					out<=225;
				end
			end
			762: begin
				if(in == 0) begin
					state<=763;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=4661;
					out<=228;
				end
				if(in == 3) begin
					state<=2761;
					out<=229;
				end
				if(in == 4) begin
					state<=6650;
					out<=230;
				end
			end
			763: begin
				if(in == 0) begin
					state<=764;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=4662;
					out<=233;
				end
				if(in == 3) begin
					state<=2762;
					out<=234;
				end
				if(in == 4) begin
					state<=6651;
					out<=235;
				end
			end
			764: begin
				if(in == 0) begin
					state<=765;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=4663;
					out<=238;
				end
				if(in == 3) begin
					state<=2763;
					out<=239;
				end
				if(in == 4) begin
					state<=6652;
					out<=240;
				end
			end
			765: begin
				if(in == 0) begin
					state<=766;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=4664;
					out<=243;
				end
				if(in == 3) begin
					state<=2764;
					out<=244;
				end
				if(in == 4) begin
					state<=6653;
					out<=245;
				end
			end
			766: begin
				if(in == 0) begin
					state<=767;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=4665;
					out<=248;
				end
				if(in == 3) begin
					state<=2765;
					out<=249;
				end
				if(in == 4) begin
					state<=6654;
					out<=250;
				end
			end
			767: begin
				if(in == 0) begin
					state<=768;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=4666;
					out<=253;
				end
				if(in == 3) begin
					state<=2766;
					out<=254;
				end
				if(in == 4) begin
					state<=6655;
					out<=255;
				end
			end
			768: begin
				if(in == 0) begin
					state<=769;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=4667;
					out<=2;
				end
				if(in == 3) begin
					state<=2767;
					out<=3;
				end
				if(in == 4) begin
					state<=6656;
					out<=4;
				end
			end
			769: begin
				if(in == 0) begin
					state<=770;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=4668;
					out<=7;
				end
				if(in == 3) begin
					state<=2768;
					out<=8;
				end
				if(in == 4) begin
					state<=6657;
					out<=9;
				end
			end
			770: begin
				if(in == 0) begin
					state<=771;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=4669;
					out<=12;
				end
				if(in == 3) begin
					state<=2769;
					out<=13;
				end
				if(in == 4) begin
					state<=6658;
					out<=14;
				end
			end
			771: begin
				if(in == 0) begin
					state<=772;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=4670;
					out<=17;
				end
				if(in == 3) begin
					state<=2770;
					out<=18;
				end
				if(in == 4) begin
					state<=6659;
					out<=19;
				end
			end
			772: begin
				if(in == 0) begin
					state<=773;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=4671;
					out<=22;
				end
				if(in == 3) begin
					state<=2771;
					out<=23;
				end
				if(in == 4) begin
					state<=6660;
					out<=24;
				end
			end
			773: begin
				if(in == 0) begin
					state<=774;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=4672;
					out<=27;
				end
				if(in == 3) begin
					state<=2772;
					out<=28;
				end
				if(in == 4) begin
					state<=6661;
					out<=29;
				end
			end
			774: begin
				if(in == 0) begin
					state<=775;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=4673;
					out<=32;
				end
				if(in == 3) begin
					state<=2773;
					out<=33;
				end
				if(in == 4) begin
					state<=6662;
					out<=34;
				end
			end
			775: begin
				if(in == 0) begin
					state<=776;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=4674;
					out<=37;
				end
				if(in == 3) begin
					state<=2774;
					out<=38;
				end
				if(in == 4) begin
					state<=6663;
					out<=39;
				end
			end
			776: begin
				if(in == 0) begin
					state<=777;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=4675;
					out<=42;
				end
				if(in == 3) begin
					state<=2775;
					out<=43;
				end
				if(in == 4) begin
					state<=6664;
					out<=44;
				end
			end
			777: begin
				if(in == 0) begin
					state<=778;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=4676;
					out<=47;
				end
				if(in == 3) begin
					state<=2776;
					out<=48;
				end
				if(in == 4) begin
					state<=6665;
					out<=49;
				end
			end
			778: begin
				if(in == 0) begin
					state<=779;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=4677;
					out<=52;
				end
				if(in == 3) begin
					state<=2777;
					out<=53;
				end
				if(in == 4) begin
					state<=6666;
					out<=54;
				end
			end
			779: begin
				if(in == 0) begin
					state<=780;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=4678;
					out<=57;
				end
				if(in == 3) begin
					state<=2778;
					out<=58;
				end
				if(in == 4) begin
					state<=6667;
					out<=59;
				end
			end
			780: begin
				if(in == 0) begin
					state<=781;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=4679;
					out<=62;
				end
				if(in == 3) begin
					state<=2779;
					out<=63;
				end
				if(in == 4) begin
					state<=6668;
					out<=64;
				end
			end
			781: begin
				if(in == 0) begin
					state<=782;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=4680;
					out<=67;
				end
				if(in == 3) begin
					state<=2780;
					out<=68;
				end
				if(in == 4) begin
					state<=6669;
					out<=69;
				end
			end
			782: begin
				if(in == 0) begin
					state<=783;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=4681;
					out<=72;
				end
				if(in == 3) begin
					state<=2781;
					out<=73;
				end
				if(in == 4) begin
					state<=6670;
					out<=74;
				end
			end
			783: begin
				if(in == 0) begin
					state<=784;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=4682;
					out<=77;
				end
				if(in == 3) begin
					state<=2782;
					out<=78;
				end
				if(in == 4) begin
					state<=6671;
					out<=79;
				end
			end
			784: begin
				if(in == 0) begin
					state<=785;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=4683;
					out<=82;
				end
				if(in == 3) begin
					state<=2783;
					out<=83;
				end
				if(in == 4) begin
					state<=6672;
					out<=84;
				end
			end
			785: begin
				if(in == 0) begin
					state<=786;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=4684;
					out<=87;
				end
				if(in == 3) begin
					state<=2784;
					out<=88;
				end
				if(in == 4) begin
					state<=6673;
					out<=89;
				end
			end
			786: begin
				if(in == 0) begin
					state<=787;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=4685;
					out<=92;
				end
				if(in == 3) begin
					state<=2785;
					out<=93;
				end
				if(in == 4) begin
					state<=6674;
					out<=94;
				end
			end
			787: begin
				if(in == 0) begin
					state<=788;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=4686;
					out<=97;
				end
				if(in == 3) begin
					state<=2786;
					out<=98;
				end
				if(in == 4) begin
					state<=6675;
					out<=99;
				end
			end
			788: begin
				if(in == 0) begin
					state<=789;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=4687;
					out<=102;
				end
				if(in == 3) begin
					state<=2787;
					out<=103;
				end
				if(in == 4) begin
					state<=6676;
					out<=104;
				end
			end
			789: begin
				if(in == 0) begin
					state<=790;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=4688;
					out<=107;
				end
				if(in == 3) begin
					state<=2788;
					out<=108;
				end
				if(in == 4) begin
					state<=6677;
					out<=109;
				end
			end
			790: begin
				if(in == 0) begin
					state<=791;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=4689;
					out<=112;
				end
				if(in == 3) begin
					state<=2789;
					out<=113;
				end
				if(in == 4) begin
					state<=6678;
					out<=114;
				end
			end
			791: begin
				if(in == 0) begin
					state<=792;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=4690;
					out<=117;
				end
				if(in == 3) begin
					state<=2790;
					out<=118;
				end
				if(in == 4) begin
					state<=6679;
					out<=119;
				end
			end
			792: begin
				if(in == 0) begin
					state<=793;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=4691;
					out<=122;
				end
				if(in == 3) begin
					state<=2791;
					out<=123;
				end
				if(in == 4) begin
					state<=6680;
					out<=124;
				end
			end
			793: begin
				if(in == 0) begin
					state<=794;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=4692;
					out<=127;
				end
				if(in == 3) begin
					state<=2792;
					out<=128;
				end
				if(in == 4) begin
					state<=6681;
					out<=129;
				end
			end
			794: begin
				if(in == 0) begin
					state<=795;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=4693;
					out<=132;
				end
				if(in == 3) begin
					state<=2793;
					out<=133;
				end
				if(in == 4) begin
					state<=6682;
					out<=134;
				end
			end
			795: begin
				if(in == 0) begin
					state<=796;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=4694;
					out<=137;
				end
				if(in == 3) begin
					state<=2794;
					out<=138;
				end
				if(in == 4) begin
					state<=6683;
					out<=139;
				end
			end
			796: begin
				if(in == 0) begin
					state<=797;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=4695;
					out<=142;
				end
				if(in == 3) begin
					state<=2795;
					out<=143;
				end
				if(in == 4) begin
					state<=6684;
					out<=144;
				end
			end
			797: begin
				if(in == 0) begin
					state<=798;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=4696;
					out<=147;
				end
				if(in == 3) begin
					state<=2796;
					out<=148;
				end
				if(in == 4) begin
					state<=6685;
					out<=149;
				end
			end
			798: begin
				if(in == 0) begin
					state<=799;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=4697;
					out<=152;
				end
				if(in == 3) begin
					state<=2797;
					out<=153;
				end
				if(in == 4) begin
					state<=6686;
					out<=154;
				end
			end
			799: begin
				if(in == 0) begin
					state<=810;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=4708;
					out<=157;
				end
				if(in == 3) begin
					state<=2808;
					out<=158;
				end
				if(in == 4) begin
					state<=6697;
					out<=159;
				end
			end
			800: begin
				if(in == 0) begin
					state<=801;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=4699;
					out<=162;
				end
				if(in == 3) begin
					state<=2799;
					out<=163;
				end
				if(in == 4) begin
					state<=6688;
					out<=164;
				end
			end
			801: begin
				if(in == 0) begin
					state<=802;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=4700;
					out<=167;
				end
				if(in == 3) begin
					state<=2800;
					out<=168;
				end
				if(in == 4) begin
					state<=6689;
					out<=169;
				end
			end
			802: begin
				if(in == 0) begin
					state<=803;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=4701;
					out<=172;
				end
				if(in == 3) begin
					state<=2801;
					out<=173;
				end
				if(in == 4) begin
					state<=6690;
					out<=174;
				end
			end
			803: begin
				if(in == 0) begin
					state<=804;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=4702;
					out<=177;
				end
				if(in == 3) begin
					state<=2802;
					out<=178;
				end
				if(in == 4) begin
					state<=6691;
					out<=179;
				end
			end
			804: begin
				if(in == 0) begin
					state<=805;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=4703;
					out<=182;
				end
				if(in == 3) begin
					state<=2803;
					out<=183;
				end
				if(in == 4) begin
					state<=6692;
					out<=184;
				end
			end
			805: begin
				if(in == 0) begin
					state<=806;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=4704;
					out<=187;
				end
				if(in == 3) begin
					state<=2804;
					out<=188;
				end
				if(in == 4) begin
					state<=6693;
					out<=189;
				end
			end
			806: begin
				if(in == 0) begin
					state<=807;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=4705;
					out<=192;
				end
				if(in == 3) begin
					state<=2805;
					out<=193;
				end
				if(in == 4) begin
					state<=6694;
					out<=194;
				end
			end
			807: begin
				if(in == 0) begin
					state<=808;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=4706;
					out<=197;
				end
				if(in == 3) begin
					state<=2806;
					out<=198;
				end
				if(in == 4) begin
					state<=6695;
					out<=199;
				end
			end
			808: begin
				if(in == 0) begin
					state<=809;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=4707;
					out<=202;
				end
				if(in == 3) begin
					state<=2807;
					out<=203;
				end
				if(in == 4) begin
					state<=6696;
					out<=204;
				end
			end
			809: begin
				if(in == 0) begin
					state<=1608;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=5497;
					out<=207;
				end
				if(in == 3) begin
					state<=3509;
					out<=208;
				end
				if(in == 4) begin
					state<=7398;
					out<=209;
				end
			end
			810: begin
				if(in == 0) begin
					state<=811;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=4709;
					out<=212;
				end
				if(in == 3) begin
					state<=2809;
					out<=213;
				end
				if(in == 4) begin
					state<=6698;
					out<=214;
				end
			end
			811: begin
				if(in == 0) begin
					state<=812;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=4710;
					out<=217;
				end
				if(in == 3) begin
					state<=2810;
					out<=218;
				end
				if(in == 4) begin
					state<=6699;
					out<=219;
				end
			end
			812: begin
				if(in == 0) begin
					state<=813;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=4711;
					out<=222;
				end
				if(in == 3) begin
					state<=2811;
					out<=223;
				end
				if(in == 4) begin
					state<=6700;
					out<=224;
				end
			end
			813: begin
				if(in == 0) begin
					state<=814;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=4712;
					out<=227;
				end
				if(in == 3) begin
					state<=2812;
					out<=228;
				end
				if(in == 4) begin
					state<=6701;
					out<=229;
				end
			end
			814: begin
				if(in == 0) begin
					state<=815;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=4713;
					out<=232;
				end
				if(in == 3) begin
					state<=2813;
					out<=233;
				end
				if(in == 4) begin
					state<=6702;
					out<=234;
				end
			end
			815: begin
				if(in == 0) begin
					state<=816;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=4714;
					out<=237;
				end
				if(in == 3) begin
					state<=2814;
					out<=238;
				end
				if(in == 4) begin
					state<=6703;
					out<=239;
				end
			end
			816: begin
				if(in == 0) begin
					state<=817;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=4715;
					out<=242;
				end
				if(in == 3) begin
					state<=2815;
					out<=243;
				end
				if(in == 4) begin
					state<=6704;
					out<=244;
				end
			end
			817: begin
				if(in == 0) begin
					state<=818;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=4716;
					out<=247;
				end
				if(in == 3) begin
					state<=2816;
					out<=248;
				end
				if(in == 4) begin
					state<=6705;
					out<=249;
				end
			end
			818: begin
				if(in == 0) begin
					state<=819;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=4717;
					out<=252;
				end
				if(in == 3) begin
					state<=2817;
					out<=253;
				end
				if(in == 4) begin
					state<=6706;
					out<=254;
				end
			end
			819: begin
				if(in == 0) begin
					state<=820;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=4718;
					out<=1;
				end
				if(in == 3) begin
					state<=2818;
					out<=2;
				end
				if(in == 4) begin
					state<=6707;
					out<=3;
				end
			end
			820: begin
				if(in == 0) begin
					state<=821;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=4719;
					out<=6;
				end
				if(in == 3) begin
					state<=2819;
					out<=7;
				end
				if(in == 4) begin
					state<=6708;
					out<=8;
				end
			end
			821: begin
				if(in == 0) begin
					state<=822;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=4720;
					out<=11;
				end
				if(in == 3) begin
					state<=2820;
					out<=12;
				end
				if(in == 4) begin
					state<=6709;
					out<=13;
				end
			end
			822: begin
				if(in == 0) begin
					state<=823;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=4721;
					out<=16;
				end
				if(in == 3) begin
					state<=2821;
					out<=17;
				end
				if(in == 4) begin
					state<=6710;
					out<=18;
				end
			end
			823: begin
				if(in == 0) begin
					state<=824;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=4722;
					out<=21;
				end
				if(in == 3) begin
					state<=2822;
					out<=22;
				end
				if(in == 4) begin
					state<=6711;
					out<=23;
				end
			end
			824: begin
				if(in == 0) begin
					state<=825;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=4723;
					out<=26;
				end
				if(in == 3) begin
					state<=2823;
					out<=27;
				end
				if(in == 4) begin
					state<=6712;
					out<=28;
				end
			end
			825: begin
				if(in == 0) begin
					state<=826;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=4724;
					out<=31;
				end
				if(in == 3) begin
					state<=2824;
					out<=32;
				end
				if(in == 4) begin
					state<=6713;
					out<=33;
				end
			end
			826: begin
				if(in == 0) begin
					state<=827;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=4725;
					out<=36;
				end
				if(in == 3) begin
					state<=2825;
					out<=37;
				end
				if(in == 4) begin
					state<=6714;
					out<=38;
				end
			end
			827: begin
				if(in == 0) begin
					state<=828;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=4726;
					out<=41;
				end
				if(in == 3) begin
					state<=2826;
					out<=42;
				end
				if(in == 4) begin
					state<=6715;
					out<=43;
				end
			end
			828: begin
				if(in == 0) begin
					state<=829;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=4727;
					out<=46;
				end
				if(in == 3) begin
					state<=2827;
					out<=47;
				end
				if(in == 4) begin
					state<=6716;
					out<=48;
				end
			end
			829: begin
				if(in == 0) begin
					state<=830;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=4728;
					out<=51;
				end
				if(in == 3) begin
					state<=2828;
					out<=52;
				end
				if(in == 4) begin
					state<=6717;
					out<=53;
				end
			end
			830: begin
				if(in == 0) begin
					state<=831;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=4729;
					out<=56;
				end
				if(in == 3) begin
					state<=2829;
					out<=57;
				end
				if(in == 4) begin
					state<=6718;
					out<=58;
				end
			end
			831: begin
				if(in == 0) begin
					state<=832;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=4730;
					out<=61;
				end
				if(in == 3) begin
					state<=2830;
					out<=62;
				end
				if(in == 4) begin
					state<=6719;
					out<=63;
				end
			end
			832: begin
				if(in == 0) begin
					state<=833;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=4731;
					out<=66;
				end
				if(in == 3) begin
					state<=2831;
					out<=67;
				end
				if(in == 4) begin
					state<=6720;
					out<=68;
				end
			end
			833: begin
				if(in == 0) begin
					state<=834;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=4732;
					out<=71;
				end
				if(in == 3) begin
					state<=2832;
					out<=72;
				end
				if(in == 4) begin
					state<=6721;
					out<=73;
				end
			end
			834: begin
				if(in == 0) begin
					state<=835;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=4733;
					out<=76;
				end
				if(in == 3) begin
					state<=2833;
					out<=77;
				end
				if(in == 4) begin
					state<=6722;
					out<=78;
				end
			end
			835: begin
				if(in == 0) begin
					state<=836;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=4734;
					out<=81;
				end
				if(in == 3) begin
					state<=2834;
					out<=82;
				end
				if(in == 4) begin
					state<=6723;
					out<=83;
				end
			end
			836: begin
				if(in == 0) begin
					state<=837;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=4735;
					out<=86;
				end
				if(in == 3) begin
					state<=2835;
					out<=87;
				end
				if(in == 4) begin
					state<=6724;
					out<=88;
				end
			end
			837: begin
				if(in == 0) begin
					state<=838;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=4736;
					out<=91;
				end
				if(in == 3) begin
					state<=2836;
					out<=92;
				end
				if(in == 4) begin
					state<=6725;
					out<=93;
				end
			end
			838: begin
				if(in == 0) begin
					state<=839;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=4737;
					out<=96;
				end
				if(in == 3) begin
					state<=2837;
					out<=97;
				end
				if(in == 4) begin
					state<=6726;
					out<=98;
				end
			end
			839: begin
				if(in == 0) begin
					state<=840;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=4738;
					out<=101;
				end
				if(in == 3) begin
					state<=2838;
					out<=102;
				end
				if(in == 4) begin
					state<=6727;
					out<=103;
				end
			end
			840: begin
				if(in == 0) begin
					state<=841;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=4739;
					out<=106;
				end
				if(in == 3) begin
					state<=2839;
					out<=107;
				end
				if(in == 4) begin
					state<=6728;
					out<=108;
				end
			end
			841: begin
				if(in == 0) begin
					state<=842;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=4740;
					out<=111;
				end
				if(in == 3) begin
					state<=2840;
					out<=112;
				end
				if(in == 4) begin
					state<=6729;
					out<=113;
				end
			end
			842: begin
				if(in == 0) begin
					state<=843;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=4741;
					out<=116;
				end
				if(in == 3) begin
					state<=2841;
					out<=117;
				end
				if(in == 4) begin
					state<=6730;
					out<=118;
				end
			end
			843: begin
				if(in == 0) begin
					state<=844;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=4742;
					out<=121;
				end
				if(in == 3) begin
					state<=2842;
					out<=122;
				end
				if(in == 4) begin
					state<=6731;
					out<=123;
				end
			end
			844: begin
				if(in == 0) begin
					state<=845;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=4743;
					out<=126;
				end
				if(in == 3) begin
					state<=2843;
					out<=127;
				end
				if(in == 4) begin
					state<=6732;
					out<=128;
				end
			end
			845: begin
				if(in == 0) begin
					state<=846;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=4744;
					out<=131;
				end
				if(in == 3) begin
					state<=2844;
					out<=132;
				end
				if(in == 4) begin
					state<=6733;
					out<=133;
				end
			end
			846: begin
				if(in == 0) begin
					state<=847;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=4745;
					out<=136;
				end
				if(in == 3) begin
					state<=2845;
					out<=137;
				end
				if(in == 4) begin
					state<=6734;
					out<=138;
				end
			end
			847: begin
				if(in == 0) begin
					state<=848;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=4746;
					out<=141;
				end
				if(in == 3) begin
					state<=2846;
					out<=142;
				end
				if(in == 4) begin
					state<=6735;
					out<=143;
				end
			end
			848: begin
				if(in == 0) begin
					state<=849;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=4747;
					out<=146;
				end
				if(in == 3) begin
					state<=2847;
					out<=147;
				end
				if(in == 4) begin
					state<=6736;
					out<=148;
				end
			end
			849: begin
				if(in == 0) begin
					state<=850;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=4748;
					out<=151;
				end
				if(in == 3) begin
					state<=2848;
					out<=152;
				end
				if(in == 4) begin
					state<=6737;
					out<=153;
				end
			end
			850: begin
				if(in == 0) begin
					state<=851;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=4749;
					out<=156;
				end
				if(in == 3) begin
					state<=2849;
					out<=157;
				end
				if(in == 4) begin
					state<=6738;
					out<=158;
				end
			end
			851: begin
				if(in == 0) begin
					state<=852;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=4750;
					out<=161;
				end
				if(in == 3) begin
					state<=2850;
					out<=162;
				end
				if(in == 4) begin
					state<=6739;
					out<=163;
				end
			end
			852: begin
				if(in == 0) begin
					state<=853;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=4751;
					out<=166;
				end
				if(in == 3) begin
					state<=2851;
					out<=167;
				end
				if(in == 4) begin
					state<=6740;
					out<=168;
				end
			end
			853: begin
				if(in == 0) begin
					state<=854;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=4752;
					out<=171;
				end
				if(in == 3) begin
					state<=2852;
					out<=172;
				end
				if(in == 4) begin
					state<=6741;
					out<=173;
				end
			end
			854: begin
				if(in == 0) begin
					state<=855;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=4753;
					out<=176;
				end
				if(in == 3) begin
					state<=2853;
					out<=177;
				end
				if(in == 4) begin
					state<=6742;
					out<=178;
				end
			end
			855: begin
				if(in == 0) begin
					state<=856;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=4754;
					out<=181;
				end
				if(in == 3) begin
					state<=2854;
					out<=182;
				end
				if(in == 4) begin
					state<=6743;
					out<=183;
				end
			end
			856: begin
				if(in == 0) begin
					state<=857;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=4755;
					out<=186;
				end
				if(in == 3) begin
					state<=2855;
					out<=187;
				end
				if(in == 4) begin
					state<=6744;
					out<=188;
				end
			end
			857: begin
				if(in == 0) begin
					state<=858;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=4756;
					out<=191;
				end
				if(in == 3) begin
					state<=2856;
					out<=192;
				end
				if(in == 4) begin
					state<=6745;
					out<=193;
				end
			end
			858: begin
				if(in == 0) begin
					state<=859;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=4757;
					out<=196;
				end
				if(in == 3) begin
					state<=2857;
					out<=197;
				end
				if(in == 4) begin
					state<=6746;
					out<=198;
				end
			end
			859: begin
				if(in == 0) begin
					state<=860;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=4758;
					out<=201;
				end
				if(in == 3) begin
					state<=2858;
					out<=202;
				end
				if(in == 4) begin
					state<=6747;
					out<=203;
				end
			end
			860: begin
				if(in == 0) begin
					state<=861;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=4759;
					out<=206;
				end
				if(in == 3) begin
					state<=2859;
					out<=207;
				end
				if(in == 4) begin
					state<=6748;
					out<=208;
				end
			end
			861: begin
				if(in == 0) begin
					state<=862;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=4760;
					out<=211;
				end
				if(in == 3) begin
					state<=2860;
					out<=212;
				end
				if(in == 4) begin
					state<=6749;
					out<=213;
				end
			end
			862: begin
				if(in == 0) begin
					state<=863;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=4761;
					out<=216;
				end
				if(in == 3) begin
					state<=2861;
					out<=217;
				end
				if(in == 4) begin
					state<=6750;
					out<=218;
				end
			end
			863: begin
				if(in == 0) begin
					state<=864;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=4762;
					out<=221;
				end
				if(in == 3) begin
					state<=2862;
					out<=222;
				end
				if(in == 4) begin
					state<=6751;
					out<=223;
				end
			end
			864: begin
				if(in == 0) begin
					state<=865;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=4763;
					out<=226;
				end
				if(in == 3) begin
					state<=2863;
					out<=227;
				end
				if(in == 4) begin
					state<=6752;
					out<=228;
				end
			end
			865: begin
				if(in == 0) begin
					state<=866;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=4764;
					out<=231;
				end
				if(in == 3) begin
					state<=2864;
					out<=232;
				end
				if(in == 4) begin
					state<=6753;
					out<=233;
				end
			end
			866: begin
				if(in == 0) begin
					state<=867;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=4765;
					out<=236;
				end
				if(in == 3) begin
					state<=2865;
					out<=237;
				end
				if(in == 4) begin
					state<=6754;
					out<=238;
				end
			end
			867: begin
				if(in == 0) begin
					state<=868;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=4766;
					out<=241;
				end
				if(in == 3) begin
					state<=2866;
					out<=242;
				end
				if(in == 4) begin
					state<=6755;
					out<=243;
				end
			end
			868: begin
				if(in == 0) begin
					state<=869;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=4767;
					out<=246;
				end
				if(in == 3) begin
					state<=2867;
					out<=247;
				end
				if(in == 4) begin
					state<=6756;
					out<=248;
				end
			end
			869: begin
				if(in == 0) begin
					state<=870;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=4768;
					out<=251;
				end
				if(in == 3) begin
					state<=2868;
					out<=252;
				end
				if(in == 4) begin
					state<=6757;
					out<=253;
				end
			end
			870: begin
				if(in == 0) begin
					state<=871;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=4769;
					out<=0;
				end
				if(in == 3) begin
					state<=2869;
					out<=1;
				end
				if(in == 4) begin
					state<=6758;
					out<=2;
				end
			end
			871: begin
				if(in == 0) begin
					state<=872;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=4770;
					out<=5;
				end
				if(in == 3) begin
					state<=2870;
					out<=6;
				end
				if(in == 4) begin
					state<=6759;
					out<=7;
				end
			end
			872: begin
				if(in == 0) begin
					state<=873;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=4771;
					out<=10;
				end
				if(in == 3) begin
					state<=2871;
					out<=11;
				end
				if(in == 4) begin
					state<=6760;
					out<=12;
				end
			end
			873: begin
				if(in == 0) begin
					state<=874;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=4772;
					out<=15;
				end
				if(in == 3) begin
					state<=2872;
					out<=16;
				end
				if(in == 4) begin
					state<=6761;
					out<=17;
				end
			end
			874: begin
				if(in == 0) begin
					state<=875;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=4773;
					out<=20;
				end
				if(in == 3) begin
					state<=2873;
					out<=21;
				end
				if(in == 4) begin
					state<=6762;
					out<=22;
				end
			end
			875: begin
				if(in == 0) begin
					state<=876;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=4774;
					out<=25;
				end
				if(in == 3) begin
					state<=2874;
					out<=26;
				end
				if(in == 4) begin
					state<=6763;
					out<=27;
				end
			end
			876: begin
				if(in == 0) begin
					state<=877;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=4775;
					out<=30;
				end
				if(in == 3) begin
					state<=2875;
					out<=31;
				end
				if(in == 4) begin
					state<=6764;
					out<=32;
				end
			end
			877: begin
				if(in == 0) begin
					state<=878;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=4776;
					out<=35;
				end
				if(in == 3) begin
					state<=2876;
					out<=36;
				end
				if(in == 4) begin
					state<=6765;
					out<=37;
				end
			end
			878: begin
				if(in == 0) begin
					state<=879;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=4777;
					out<=40;
				end
				if(in == 3) begin
					state<=2877;
					out<=41;
				end
				if(in == 4) begin
					state<=6766;
					out<=42;
				end
			end
			879: begin
				if(in == 0) begin
					state<=880;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=4778;
					out<=45;
				end
				if(in == 3) begin
					state<=2878;
					out<=46;
				end
				if(in == 4) begin
					state<=6767;
					out<=47;
				end
			end
			880: begin
				if(in == 0) begin
					state<=881;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=4779;
					out<=50;
				end
				if(in == 3) begin
					state<=2879;
					out<=51;
				end
				if(in == 4) begin
					state<=6768;
					out<=52;
				end
			end
			881: begin
				if(in == 0) begin
					state<=882;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=4780;
					out<=55;
				end
				if(in == 3) begin
					state<=2880;
					out<=56;
				end
				if(in == 4) begin
					state<=6769;
					out<=57;
				end
			end
			882: begin
				if(in == 0) begin
					state<=883;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=4781;
					out<=60;
				end
				if(in == 3) begin
					state<=2881;
					out<=61;
				end
				if(in == 4) begin
					state<=6770;
					out<=62;
				end
			end
			883: begin
				if(in == 0) begin
					state<=884;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=4782;
					out<=65;
				end
				if(in == 3) begin
					state<=2882;
					out<=66;
				end
				if(in == 4) begin
					state<=6771;
					out<=67;
				end
			end
			884: begin
				if(in == 0) begin
					state<=885;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=4783;
					out<=70;
				end
				if(in == 3) begin
					state<=2883;
					out<=71;
				end
				if(in == 4) begin
					state<=6772;
					out<=72;
				end
			end
			885: begin
				if(in == 0) begin
					state<=886;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=4784;
					out<=75;
				end
				if(in == 3) begin
					state<=2884;
					out<=76;
				end
				if(in == 4) begin
					state<=6773;
					out<=77;
				end
			end
			886: begin
				if(in == 0) begin
					state<=887;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=4785;
					out<=80;
				end
				if(in == 3) begin
					state<=2885;
					out<=81;
				end
				if(in == 4) begin
					state<=6774;
					out<=82;
				end
			end
			887: begin
				if(in == 0) begin
					state<=888;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=4786;
					out<=85;
				end
				if(in == 3) begin
					state<=2886;
					out<=86;
				end
				if(in == 4) begin
					state<=6775;
					out<=87;
				end
			end
			888: begin
				if(in == 0) begin
					state<=889;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=4787;
					out<=90;
				end
				if(in == 3) begin
					state<=2887;
					out<=91;
				end
				if(in == 4) begin
					state<=6776;
					out<=92;
				end
			end
			889: begin
				if(in == 0) begin
					state<=890;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=4788;
					out<=95;
				end
				if(in == 3) begin
					state<=2888;
					out<=96;
				end
				if(in == 4) begin
					state<=6777;
					out<=97;
				end
			end
			890: begin
				if(in == 0) begin
					state<=891;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=4789;
					out<=100;
				end
				if(in == 3) begin
					state<=2889;
					out<=101;
				end
				if(in == 4) begin
					state<=6778;
					out<=102;
				end
			end
			891: begin
				if(in == 0) begin
					state<=892;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=4790;
					out<=105;
				end
				if(in == 3) begin
					state<=2890;
					out<=106;
				end
				if(in == 4) begin
					state<=6779;
					out<=107;
				end
			end
			892: begin
				if(in == 0) begin
					state<=893;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=4791;
					out<=110;
				end
				if(in == 3) begin
					state<=2891;
					out<=111;
				end
				if(in == 4) begin
					state<=6780;
					out<=112;
				end
			end
			893: begin
				if(in == 0) begin
					state<=894;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=4792;
					out<=115;
				end
				if(in == 3) begin
					state<=2892;
					out<=116;
				end
				if(in == 4) begin
					state<=6781;
					out<=117;
				end
			end
			894: begin
				if(in == 0) begin
					state<=895;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=4793;
					out<=120;
				end
				if(in == 3) begin
					state<=2893;
					out<=121;
				end
				if(in == 4) begin
					state<=6782;
					out<=122;
				end
			end
			895: begin
				if(in == 0) begin
					state<=896;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=4794;
					out<=125;
				end
				if(in == 3) begin
					state<=2894;
					out<=126;
				end
				if(in == 4) begin
					state<=6783;
					out<=127;
				end
			end
			896: begin
				if(in == 0) begin
					state<=897;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=4795;
					out<=130;
				end
				if(in == 3) begin
					state<=2895;
					out<=131;
				end
				if(in == 4) begin
					state<=6784;
					out<=132;
				end
			end
			897: begin
				if(in == 0) begin
					state<=898;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=4796;
					out<=135;
				end
				if(in == 3) begin
					state<=2896;
					out<=136;
				end
				if(in == 4) begin
					state<=6785;
					out<=137;
				end
			end
			898: begin
				if(in == 0) begin
					state<=899;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=4797;
					out<=140;
				end
				if(in == 3) begin
					state<=2897;
					out<=141;
				end
				if(in == 4) begin
					state<=6786;
					out<=142;
				end
			end
			899: begin
				if(in == 0) begin
					state<=800;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=4698;
					out<=145;
				end
				if(in == 3) begin
					state<=2798;
					out<=146;
				end
				if(in == 4) begin
					state<=6687;
					out<=147;
				end
			end
			900: begin
				if(in == 0) begin
					state<=901;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=4799;
					out<=150;
				end
				if(in == 3) begin
					state<=2277;
					out<=151;
				end
				if(in == 4) begin
					state<=6166;
					out<=152;
				end
			end
			901: begin
				if(in == 0) begin
					state<=902;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=4800;
					out<=155;
				end
				if(in == 3) begin
					state<=2278;
					out<=156;
				end
				if(in == 4) begin
					state<=6167;
					out<=157;
				end
			end
			902: begin
				if(in == 0) begin
					state<=903;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=4801;
					out<=160;
				end
				if(in == 3) begin
					state<=2279;
					out<=161;
				end
				if(in == 4) begin
					state<=6168;
					out<=162;
				end
			end
			903: begin
				if(in == 0) begin
					state<=904;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=4802;
					out<=165;
				end
				if(in == 3) begin
					state<=2280;
					out<=166;
				end
				if(in == 4) begin
					state<=6169;
					out<=167;
				end
			end
			904: begin
				if(in == 0) begin
					state<=905;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=4803;
					out<=170;
				end
				if(in == 3) begin
					state<=2281;
					out<=171;
				end
				if(in == 4) begin
					state<=6170;
					out<=172;
				end
			end
			905: begin
				if(in == 0) begin
					state<=906;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=4804;
					out<=175;
				end
				if(in == 3) begin
					state<=2282;
					out<=176;
				end
				if(in == 4) begin
					state<=6171;
					out<=177;
				end
			end
			906: begin
				if(in == 0) begin
					state<=907;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=4805;
					out<=180;
				end
				if(in == 3) begin
					state<=2283;
					out<=181;
				end
				if(in == 4) begin
					state<=6172;
					out<=182;
				end
			end
			907: begin
				if(in == 0) begin
					state<=908;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=4806;
					out<=185;
				end
				if(in == 3) begin
					state<=2284;
					out<=186;
				end
				if(in == 4) begin
					state<=6173;
					out<=187;
				end
			end
			908: begin
				if(in == 0) begin
					state<=909;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=4807;
					out<=190;
				end
				if(in == 3) begin
					state<=2285;
					out<=191;
				end
				if(in == 4) begin
					state<=6174;
					out<=192;
				end
			end
			909: begin
				if(in == 0) begin
					state<=910;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=4808;
					out<=195;
				end
				if(in == 3) begin
					state<=2286;
					out<=196;
				end
				if(in == 4) begin
					state<=6175;
					out<=197;
				end
			end
			910: begin
				if(in == 0) begin
					state<=911;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=4809;
					out<=200;
				end
				if(in == 3) begin
					state<=2287;
					out<=201;
				end
				if(in == 4) begin
					state<=6176;
					out<=202;
				end
			end
			911: begin
				if(in == 0) begin
					state<=912;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=4810;
					out<=205;
				end
				if(in == 3) begin
					state<=2288;
					out<=206;
				end
				if(in == 4) begin
					state<=6177;
					out<=207;
				end
			end
			912: begin
				if(in == 0) begin
					state<=913;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=4811;
					out<=210;
				end
				if(in == 3) begin
					state<=2289;
					out<=211;
				end
				if(in == 4) begin
					state<=6178;
					out<=212;
				end
			end
			913: begin
				if(in == 0) begin
					state<=914;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=4812;
					out<=215;
				end
				if(in == 3) begin
					state<=2290;
					out<=216;
				end
				if(in == 4) begin
					state<=6179;
					out<=217;
				end
			end
			914: begin
				if(in == 0) begin
					state<=915;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=4813;
					out<=220;
				end
				if(in == 3) begin
					state<=2291;
					out<=221;
				end
				if(in == 4) begin
					state<=6180;
					out<=222;
				end
			end
			915: begin
				if(in == 0) begin
					state<=916;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=4814;
					out<=225;
				end
				if(in == 3) begin
					state<=2292;
					out<=226;
				end
				if(in == 4) begin
					state<=6181;
					out<=227;
				end
			end
			916: begin
				if(in == 0) begin
					state<=917;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=4815;
					out<=230;
				end
				if(in == 3) begin
					state<=2293;
					out<=231;
				end
				if(in == 4) begin
					state<=6182;
					out<=232;
				end
			end
			917: begin
				if(in == 0) begin
					state<=918;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=4816;
					out<=235;
				end
				if(in == 3) begin
					state<=2294;
					out<=236;
				end
				if(in == 4) begin
					state<=6183;
					out<=237;
				end
			end
			918: begin
				if(in == 0) begin
					state<=919;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=4817;
					out<=240;
				end
				if(in == 3) begin
					state<=2295;
					out<=241;
				end
				if(in == 4) begin
					state<=6184;
					out<=242;
				end
			end
			919: begin
				if(in == 0) begin
					state<=920;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=4818;
					out<=245;
				end
				if(in == 3) begin
					state<=2296;
					out<=246;
				end
				if(in == 4) begin
					state<=6185;
					out<=247;
				end
			end
			920: begin
				if(in == 0) begin
					state<=921;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=4819;
					out<=250;
				end
				if(in == 3) begin
					state<=2297;
					out<=251;
				end
				if(in == 4) begin
					state<=6186;
					out<=252;
				end
			end
			921: begin
				if(in == 0) begin
					state<=922;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=4820;
					out<=255;
				end
				if(in == 3) begin
					state<=2298;
					out<=0;
				end
				if(in == 4) begin
					state<=6187;
					out<=1;
				end
			end
			922: begin
				if(in == 0) begin
					state<=923;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=4821;
					out<=4;
				end
				if(in == 3) begin
					state<=2299;
					out<=5;
				end
				if(in == 4) begin
					state<=6188;
					out<=6;
				end
			end
			923: begin
				if(in == 0) begin
					state<=924;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=4822;
					out<=9;
				end
				if(in == 3) begin
					state<=2300;
					out<=10;
				end
				if(in == 4) begin
					state<=6189;
					out<=11;
				end
			end
			924: begin
				if(in == 0) begin
					state<=925;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=4823;
					out<=14;
				end
				if(in == 3) begin
					state<=2301;
					out<=15;
				end
				if(in == 4) begin
					state<=6190;
					out<=16;
				end
			end
			925: begin
				if(in == 0) begin
					state<=926;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=4824;
					out<=19;
				end
				if(in == 3) begin
					state<=2302;
					out<=20;
				end
				if(in == 4) begin
					state<=6191;
					out<=21;
				end
			end
			926: begin
				if(in == 0) begin
					state<=927;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=4825;
					out<=24;
				end
				if(in == 3) begin
					state<=2303;
					out<=25;
				end
				if(in == 4) begin
					state<=6192;
					out<=26;
				end
			end
			927: begin
				if(in == 0) begin
					state<=928;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=4826;
					out<=29;
				end
				if(in == 3) begin
					state<=2304;
					out<=30;
				end
				if(in == 4) begin
					state<=6193;
					out<=31;
				end
			end
			928: begin
				if(in == 0) begin
					state<=929;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=4827;
					out<=34;
				end
				if(in == 3) begin
					state<=2305;
					out<=35;
				end
				if(in == 4) begin
					state<=6194;
					out<=36;
				end
			end
			929: begin
				if(in == 0) begin
					state<=930;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=4828;
					out<=39;
				end
				if(in == 3) begin
					state<=2306;
					out<=40;
				end
				if(in == 4) begin
					state<=6195;
					out<=41;
				end
			end
			930: begin
				if(in == 0) begin
					state<=931;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=4829;
					out<=44;
				end
				if(in == 3) begin
					state<=2307;
					out<=45;
				end
				if(in == 4) begin
					state<=6196;
					out<=46;
				end
			end
			931: begin
				if(in == 0) begin
					state<=932;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=4830;
					out<=49;
				end
				if(in == 3) begin
					state<=2308;
					out<=50;
				end
				if(in == 4) begin
					state<=6197;
					out<=51;
				end
			end
			932: begin
				if(in == 0) begin
					state<=933;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=4831;
					out<=54;
				end
				if(in == 3) begin
					state<=2309;
					out<=55;
				end
				if(in == 4) begin
					state<=6198;
					out<=56;
				end
			end
			933: begin
				if(in == 0) begin
					state<=934;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=4832;
					out<=59;
				end
				if(in == 3) begin
					state<=2310;
					out<=60;
				end
				if(in == 4) begin
					state<=6199;
					out<=61;
				end
			end
			934: begin
				if(in == 0) begin
					state<=935;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=4833;
					out<=64;
				end
				if(in == 3) begin
					state<=2311;
					out<=65;
				end
				if(in == 4) begin
					state<=6200;
					out<=66;
				end
			end
			935: begin
				if(in == 0) begin
					state<=936;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=4834;
					out<=69;
				end
				if(in == 3) begin
					state<=2312;
					out<=70;
				end
				if(in == 4) begin
					state<=6201;
					out<=71;
				end
			end
			936: begin
				if(in == 0) begin
					state<=937;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=4835;
					out<=74;
				end
				if(in == 3) begin
					state<=2313;
					out<=75;
				end
				if(in == 4) begin
					state<=6202;
					out<=76;
				end
			end
			937: begin
				if(in == 0) begin
					state<=938;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=4836;
					out<=79;
				end
				if(in == 3) begin
					state<=2314;
					out<=80;
				end
				if(in == 4) begin
					state<=6203;
					out<=81;
				end
			end
			938: begin
				if(in == 0) begin
					state<=939;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=4837;
					out<=84;
				end
				if(in == 3) begin
					state<=2315;
					out<=85;
				end
				if(in == 4) begin
					state<=6204;
					out<=86;
				end
			end
			939: begin
				if(in == 0) begin
					state<=940;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=4838;
					out<=89;
				end
				if(in == 3) begin
					state<=2316;
					out<=90;
				end
				if(in == 4) begin
					state<=6205;
					out<=91;
				end
			end
			940: begin
				if(in == 0) begin
					state<=941;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=4839;
					out<=94;
				end
				if(in == 3) begin
					state<=2317;
					out<=95;
				end
				if(in == 4) begin
					state<=6206;
					out<=96;
				end
			end
			941: begin
				if(in == 0) begin
					state<=942;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=4840;
					out<=99;
				end
				if(in == 3) begin
					state<=2318;
					out<=100;
				end
				if(in == 4) begin
					state<=6207;
					out<=101;
				end
			end
			942: begin
				if(in == 0) begin
					state<=943;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=4841;
					out<=104;
				end
				if(in == 3) begin
					state<=2319;
					out<=105;
				end
				if(in == 4) begin
					state<=6208;
					out<=106;
				end
			end
			943: begin
				if(in == 0) begin
					state<=944;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=4842;
					out<=109;
				end
				if(in == 3) begin
					state<=2320;
					out<=110;
				end
				if(in == 4) begin
					state<=6209;
					out<=111;
				end
			end
			944: begin
				if(in == 0) begin
					state<=945;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=4843;
					out<=114;
				end
				if(in == 3) begin
					state<=2321;
					out<=115;
				end
				if(in == 4) begin
					state<=6210;
					out<=116;
				end
			end
			945: begin
				if(in == 0) begin
					state<=946;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=4844;
					out<=119;
				end
				if(in == 3) begin
					state<=2322;
					out<=120;
				end
				if(in == 4) begin
					state<=6211;
					out<=121;
				end
			end
			946: begin
				if(in == 0) begin
					state<=947;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=4845;
					out<=124;
				end
				if(in == 3) begin
					state<=2323;
					out<=125;
				end
				if(in == 4) begin
					state<=6212;
					out<=126;
				end
			end
			947: begin
				if(in == 0) begin
					state<=948;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=4846;
					out<=129;
				end
				if(in == 3) begin
					state<=2324;
					out<=130;
				end
				if(in == 4) begin
					state<=6213;
					out<=131;
				end
			end
			948: begin
				if(in == 0) begin
					state<=949;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=4847;
					out<=134;
				end
				if(in == 3) begin
					state<=2898;
					out<=135;
				end
				if(in == 4) begin
					state<=6787;
					out<=136;
				end
			end
			949: begin
				if(in == 0) begin
					state<=950;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=4848;
					out<=139;
				end
				if(in == 3) begin
					state<=2899;
					out<=140;
				end
				if(in == 4) begin
					state<=6788;
					out<=141;
				end
			end
			950: begin
				if(in == 0) begin
					state<=951;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=4849;
					out<=144;
				end
				if(in == 3) begin
					state<=2900;
					out<=145;
				end
				if(in == 4) begin
					state<=6789;
					out<=146;
				end
			end
			951: begin
				if(in == 0) begin
					state<=952;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=4850;
					out<=149;
				end
				if(in == 3) begin
					state<=2901;
					out<=150;
				end
				if(in == 4) begin
					state<=6790;
					out<=151;
				end
			end
			952: begin
				if(in == 0) begin
					state<=953;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=4851;
					out<=154;
				end
				if(in == 3) begin
					state<=2902;
					out<=155;
				end
				if(in == 4) begin
					state<=6791;
					out<=156;
				end
			end
			953: begin
				if(in == 0) begin
					state<=954;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=4852;
					out<=159;
				end
				if(in == 3) begin
					state<=2903;
					out<=160;
				end
				if(in == 4) begin
					state<=6792;
					out<=161;
				end
			end
			954: begin
				if(in == 0) begin
					state<=955;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=4853;
					out<=164;
				end
				if(in == 3) begin
					state<=2904;
					out<=165;
				end
				if(in == 4) begin
					state<=6793;
					out<=166;
				end
			end
			955: begin
				if(in == 0) begin
					state<=956;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=4854;
					out<=169;
				end
				if(in == 3) begin
					state<=2905;
					out<=170;
				end
				if(in == 4) begin
					state<=6794;
					out<=171;
				end
			end
			956: begin
				if(in == 0) begin
					state<=957;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=4855;
					out<=174;
				end
				if(in == 3) begin
					state<=2906;
					out<=175;
				end
				if(in == 4) begin
					state<=6795;
					out<=176;
				end
			end
			957: begin
				if(in == 0) begin
					state<=958;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=4856;
					out<=179;
				end
				if(in == 3) begin
					state<=2907;
					out<=180;
				end
				if(in == 4) begin
					state<=6796;
					out<=181;
				end
			end
			958: begin
				if(in == 0) begin
					state<=959;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=4857;
					out<=184;
				end
				if(in == 3) begin
					state<=2908;
					out<=185;
				end
				if(in == 4) begin
					state<=6797;
					out<=186;
				end
			end
			959: begin
				if(in == 0) begin
					state<=960;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=4858;
					out<=189;
				end
				if(in == 3) begin
					state<=2909;
					out<=190;
				end
				if(in == 4) begin
					state<=6798;
					out<=191;
				end
			end
			960: begin
				if(in == 0) begin
					state<=961;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=4859;
					out<=194;
				end
				if(in == 3) begin
					state<=2910;
					out<=195;
				end
				if(in == 4) begin
					state<=6799;
					out<=196;
				end
			end
			961: begin
				if(in == 0) begin
					state<=962;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=4860;
					out<=199;
				end
				if(in == 3) begin
					state<=2911;
					out<=200;
				end
				if(in == 4) begin
					state<=6800;
					out<=201;
				end
			end
			962: begin
				if(in == 0) begin
					state<=963;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=4861;
					out<=204;
				end
				if(in == 3) begin
					state<=2912;
					out<=205;
				end
				if(in == 4) begin
					state<=6801;
					out<=206;
				end
			end
			963: begin
				if(in == 0) begin
					state<=964;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=4862;
					out<=209;
				end
				if(in == 3) begin
					state<=2913;
					out<=210;
				end
				if(in == 4) begin
					state<=6802;
					out<=211;
				end
			end
			964: begin
				if(in == 0) begin
					state<=965;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=4863;
					out<=214;
				end
				if(in == 3) begin
					state<=2914;
					out<=215;
				end
				if(in == 4) begin
					state<=6803;
					out<=216;
				end
			end
			965: begin
				if(in == 0) begin
					state<=966;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=4864;
					out<=219;
				end
				if(in == 3) begin
					state<=2915;
					out<=220;
				end
				if(in == 4) begin
					state<=6804;
					out<=221;
				end
			end
			966: begin
				if(in == 0) begin
					state<=967;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=4865;
					out<=224;
				end
				if(in == 3) begin
					state<=2916;
					out<=225;
				end
				if(in == 4) begin
					state<=6805;
					out<=226;
				end
			end
			967: begin
				if(in == 0) begin
					state<=968;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=4866;
					out<=229;
				end
				if(in == 3) begin
					state<=2917;
					out<=230;
				end
				if(in == 4) begin
					state<=6806;
					out<=231;
				end
			end
			968: begin
				if(in == 0) begin
					state<=969;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=4867;
					out<=234;
				end
				if(in == 3) begin
					state<=2918;
					out<=235;
				end
				if(in == 4) begin
					state<=6807;
					out<=236;
				end
			end
			969: begin
				if(in == 0) begin
					state<=970;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=4868;
					out<=239;
				end
				if(in == 3) begin
					state<=2919;
					out<=240;
				end
				if(in == 4) begin
					state<=6808;
					out<=241;
				end
			end
			970: begin
				if(in == 0) begin
					state<=971;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=4869;
					out<=244;
				end
				if(in == 3) begin
					state<=2920;
					out<=245;
				end
				if(in == 4) begin
					state<=6809;
					out<=246;
				end
			end
			971: begin
				if(in == 0) begin
					state<=972;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=4870;
					out<=249;
				end
				if(in == 3) begin
					state<=2921;
					out<=250;
				end
				if(in == 4) begin
					state<=6810;
					out<=251;
				end
			end
			972: begin
				if(in == 0) begin
					state<=973;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=4871;
					out<=254;
				end
				if(in == 3) begin
					state<=2922;
					out<=255;
				end
				if(in == 4) begin
					state<=6811;
					out<=0;
				end
			end
			973: begin
				if(in == 0) begin
					state<=974;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=4872;
					out<=3;
				end
				if(in == 3) begin
					state<=2923;
					out<=4;
				end
				if(in == 4) begin
					state<=6812;
					out<=5;
				end
			end
			974: begin
				if(in == 0) begin
					state<=975;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=4873;
					out<=8;
				end
				if(in == 3) begin
					state<=2924;
					out<=9;
				end
				if(in == 4) begin
					state<=6813;
					out<=10;
				end
			end
			975: begin
				if(in == 0) begin
					state<=976;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=4874;
					out<=13;
				end
				if(in == 3) begin
					state<=2925;
					out<=14;
				end
				if(in == 4) begin
					state<=6814;
					out<=15;
				end
			end
			976: begin
				if(in == 0) begin
					state<=977;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=4875;
					out<=18;
				end
				if(in == 3) begin
					state<=2926;
					out<=19;
				end
				if(in == 4) begin
					state<=6815;
					out<=20;
				end
			end
			977: begin
				if(in == 0) begin
					state<=978;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=4876;
					out<=23;
				end
				if(in == 3) begin
					state<=2927;
					out<=24;
				end
				if(in == 4) begin
					state<=6816;
					out<=25;
				end
			end
			978: begin
				if(in == 0) begin
					state<=979;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=4877;
					out<=28;
				end
				if(in == 3) begin
					state<=2928;
					out<=29;
				end
				if(in == 4) begin
					state<=6817;
					out<=30;
				end
			end
			979: begin
				if(in == 0) begin
					state<=980;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=4878;
					out<=33;
				end
				if(in == 3) begin
					state<=2325;
					out<=34;
				end
				if(in == 4) begin
					state<=6214;
					out<=35;
				end
			end
			980: begin
				if(in == 0) begin
					state<=981;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=4879;
					out<=38;
				end
				if(in == 3) begin
					state<=2326;
					out<=39;
				end
				if(in == 4) begin
					state<=6215;
					out<=40;
				end
			end
			981: begin
				if(in == 0) begin
					state<=982;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=4880;
					out<=43;
				end
				if(in == 3) begin
					state<=2327;
					out<=44;
				end
				if(in == 4) begin
					state<=6216;
					out<=45;
				end
			end
			982: begin
				if(in == 0) begin
					state<=983;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=4881;
					out<=48;
				end
				if(in == 3) begin
					state<=2328;
					out<=49;
				end
				if(in == 4) begin
					state<=6217;
					out<=50;
				end
			end
			983: begin
				if(in == 0) begin
					state<=984;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=4882;
					out<=53;
				end
				if(in == 3) begin
					state<=2329;
					out<=54;
				end
				if(in == 4) begin
					state<=6218;
					out<=55;
				end
			end
			984: begin
				if(in == 0) begin
					state<=985;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=4883;
					out<=58;
				end
				if(in == 3) begin
					state<=2330;
					out<=59;
				end
				if(in == 4) begin
					state<=6219;
					out<=60;
				end
			end
			985: begin
				if(in == 0) begin
					state<=986;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=4884;
					out<=63;
				end
				if(in == 3) begin
					state<=2331;
					out<=64;
				end
				if(in == 4) begin
					state<=6220;
					out<=65;
				end
			end
			986: begin
				if(in == 0) begin
					state<=987;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=4885;
					out<=68;
				end
				if(in == 3) begin
					state<=2332;
					out<=69;
				end
				if(in == 4) begin
					state<=6221;
					out<=70;
				end
			end
			987: begin
				if(in == 0) begin
					state<=988;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=4886;
					out<=73;
				end
				if(in == 3) begin
					state<=2333;
					out<=74;
				end
				if(in == 4) begin
					state<=6222;
					out<=75;
				end
			end
			988: begin
				if(in == 0) begin
					state<=989;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=4887;
					out<=78;
				end
				if(in == 3) begin
					state<=2334;
					out<=79;
				end
				if(in == 4) begin
					state<=6223;
					out<=80;
				end
			end
			989: begin
				if(in == 0) begin
					state<=990;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=4888;
					out<=83;
				end
				if(in == 3) begin
					state<=2335;
					out<=84;
				end
				if(in == 4) begin
					state<=6224;
					out<=85;
				end
			end
			990: begin
				if(in == 0) begin
					state<=991;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=4889;
					out<=88;
				end
				if(in == 3) begin
					state<=2336;
					out<=89;
				end
				if(in == 4) begin
					state<=6225;
					out<=90;
				end
			end
			991: begin
				if(in == 0) begin
					state<=992;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=4890;
					out<=93;
				end
				if(in == 3) begin
					state<=2337;
					out<=94;
				end
				if(in == 4) begin
					state<=6226;
					out<=95;
				end
			end
			992: begin
				if(in == 0) begin
					state<=993;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=4891;
					out<=98;
				end
				if(in == 3) begin
					state<=2338;
					out<=99;
				end
				if(in == 4) begin
					state<=6227;
					out<=100;
				end
			end
			993: begin
				if(in == 0) begin
					state<=994;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=4892;
					out<=103;
				end
				if(in == 3) begin
					state<=2339;
					out<=104;
				end
				if(in == 4) begin
					state<=6228;
					out<=105;
				end
			end
			994: begin
				if(in == 0) begin
					state<=995;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=4893;
					out<=108;
				end
				if(in == 3) begin
					state<=2340;
					out<=109;
				end
				if(in == 4) begin
					state<=6229;
					out<=110;
				end
			end
			995: begin
				if(in == 0) begin
					state<=996;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=4894;
					out<=113;
				end
				if(in == 3) begin
					state<=2341;
					out<=114;
				end
				if(in == 4) begin
					state<=6230;
					out<=115;
				end
			end
			996: begin
				if(in == 0) begin
					state<=997;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=4895;
					out<=118;
				end
				if(in == 3) begin
					state<=2342;
					out<=119;
				end
				if(in == 4) begin
					state<=6231;
					out<=120;
				end
			end
			997: begin
				if(in == 0) begin
					state<=998;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=4896;
					out<=123;
				end
				if(in == 3) begin
					state<=2343;
					out<=124;
				end
				if(in == 4) begin
					state<=6232;
					out<=125;
				end
			end
			998: begin
				if(in == 0) begin
					state<=346;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=4244;
					out<=128;
				end
				if(in == 3) begin
					state<=2929;
					out<=129;
				end
				if(in == 4) begin
					state<=6818;
					out<=130;
				end
			end
			999: begin
				if(in == 0) begin
					state<=1000;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=4898;
					out<=133;
				end
				if(in == 3) begin
					state<=2980;
					out<=134;
				end
				if(in == 4) begin
					state<=6869;
					out<=135;
				end
			end
			1000: begin
				if(in == 0) begin
					state<=1001;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=4899;
					out<=138;
				end
				if(in == 3) begin
					state<=2981;
					out<=139;
				end
				if(in == 4) begin
					state<=6870;
					out<=140;
				end
			end
			1001: begin
				if(in == 0) begin
					state<=1002;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=4900;
					out<=143;
				end
				if(in == 3) begin
					state<=2982;
					out<=144;
				end
				if(in == 4) begin
					state<=6871;
					out<=145;
				end
			end
			1002: begin
				if(in == 0) begin
					state<=1003;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=4901;
					out<=148;
				end
				if(in == 3) begin
					state<=2983;
					out<=149;
				end
				if(in == 4) begin
					state<=6872;
					out<=150;
				end
			end
			1003: begin
				if(in == 0) begin
					state<=1004;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=4902;
					out<=153;
				end
				if(in == 3) begin
					state<=2984;
					out<=154;
				end
				if(in == 4) begin
					state<=6873;
					out<=155;
				end
			end
			1004: begin
				if(in == 0) begin
					state<=1005;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=4903;
					out<=158;
				end
				if(in == 3) begin
					state<=2985;
					out<=159;
				end
				if(in == 4) begin
					state<=6874;
					out<=160;
				end
			end
			1005: begin
				if(in == 0) begin
					state<=1006;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=4904;
					out<=163;
				end
				if(in == 3) begin
					state<=2986;
					out<=164;
				end
				if(in == 4) begin
					state<=6875;
					out<=165;
				end
			end
			1006: begin
				if(in == 0) begin
					state<=1007;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=4905;
					out<=168;
				end
				if(in == 3) begin
					state<=2987;
					out<=169;
				end
				if(in == 4) begin
					state<=6876;
					out<=170;
				end
			end
			1007: begin
				if(in == 0) begin
					state<=1008;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=4906;
					out<=173;
				end
				if(in == 3) begin
					state<=2988;
					out<=174;
				end
				if(in == 4) begin
					state<=6877;
					out<=175;
				end
			end
			1008: begin
				if(in == 0) begin
					state<=1009;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=4907;
					out<=178;
				end
				if(in == 3) begin
					state<=2989;
					out<=179;
				end
				if(in == 4) begin
					state<=6878;
					out<=180;
				end
			end
			1009: begin
				if(in == 0) begin
					state<=1010;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=4908;
					out<=183;
				end
				if(in == 3) begin
					state<=2990;
					out<=184;
				end
				if(in == 4) begin
					state<=6879;
					out<=185;
				end
			end
			1010: begin
				if(in == 0) begin
					state<=1011;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=4909;
					out<=188;
				end
				if(in == 3) begin
					state<=2991;
					out<=189;
				end
				if(in == 4) begin
					state<=6880;
					out<=190;
				end
			end
			1011: begin
				if(in == 0) begin
					state<=1012;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=4910;
					out<=193;
				end
				if(in == 3) begin
					state<=2992;
					out<=194;
				end
				if(in == 4) begin
					state<=6881;
					out<=195;
				end
			end
			1012: begin
				if(in == 0) begin
					state<=1013;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=4911;
					out<=198;
				end
				if(in == 3) begin
					state<=2993;
					out<=199;
				end
				if(in == 4) begin
					state<=6882;
					out<=200;
				end
			end
			1013: begin
				if(in == 0) begin
					state<=1014;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=4912;
					out<=203;
				end
				if(in == 3) begin
					state<=2994;
					out<=204;
				end
				if(in == 4) begin
					state<=6883;
					out<=205;
				end
			end
			1014: begin
				if(in == 0) begin
					state<=1015;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=4913;
					out<=208;
				end
				if(in == 3) begin
					state<=2995;
					out<=209;
				end
				if(in == 4) begin
					state<=6884;
					out<=210;
				end
			end
			1015: begin
				if(in == 0) begin
					state<=1016;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=4914;
					out<=213;
				end
				if(in == 3) begin
					state<=2996;
					out<=214;
				end
				if(in == 4) begin
					state<=6885;
					out<=215;
				end
			end
			1016: begin
				if(in == 0) begin
					state<=1017;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=4915;
					out<=218;
				end
				if(in == 3) begin
					state<=2997;
					out<=219;
				end
				if(in == 4) begin
					state<=6886;
					out<=220;
				end
			end
			1017: begin
				if(in == 0) begin
					state<=1018;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=4916;
					out<=223;
				end
				if(in == 3) begin
					state<=2998;
					out<=224;
				end
				if(in == 4) begin
					state<=6887;
					out<=225;
				end
			end
			1018: begin
				if(in == 0) begin
					state<=1019;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=4917;
					out<=228;
				end
				if(in == 3) begin
					state<=2999;
					out<=229;
				end
				if(in == 4) begin
					state<=6888;
					out<=230;
				end
			end
			1019: begin
				if(in == 0) begin
					state<=1020;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=4918;
					out<=233;
				end
				if(in == 3) begin
					state<=3000;
					out<=234;
				end
				if(in == 4) begin
					state<=6889;
					out<=235;
				end
			end
			1020: begin
				if(in == 0) begin
					state<=1021;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=4919;
					out<=238;
				end
				if(in == 3) begin
					state<=3001;
					out<=239;
				end
				if(in == 4) begin
					state<=6890;
					out<=240;
				end
			end
			1021: begin
				if(in == 0) begin
					state<=1022;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=4920;
					out<=243;
				end
				if(in == 3) begin
					state<=3002;
					out<=244;
				end
				if(in == 4) begin
					state<=6891;
					out<=245;
				end
			end
			1022: begin
				if(in == 0) begin
					state<=1023;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=4921;
					out<=248;
				end
				if(in == 3) begin
					state<=3003;
					out<=249;
				end
				if(in == 4) begin
					state<=6892;
					out<=250;
				end
			end
			1023: begin
				if(in == 0) begin
					state<=1024;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=4922;
					out<=253;
				end
				if(in == 3) begin
					state<=3004;
					out<=254;
				end
				if(in == 4) begin
					state<=6893;
					out<=255;
				end
			end
			1024: begin
				if(in == 0) begin
					state<=1025;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=4923;
					out<=2;
				end
				if(in == 3) begin
					state<=3005;
					out<=3;
				end
				if(in == 4) begin
					state<=6894;
					out<=4;
				end
			end
			1025: begin
				if(in == 0) begin
					state<=1026;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=4924;
					out<=7;
				end
				if(in == 3) begin
					state<=3006;
					out<=8;
				end
				if(in == 4) begin
					state<=6895;
					out<=9;
				end
			end
			1026: begin
				if(in == 0) begin
					state<=1027;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=4925;
					out<=12;
				end
				if(in == 3) begin
					state<=3007;
					out<=13;
				end
				if(in == 4) begin
					state<=6896;
					out<=14;
				end
			end
			1027: begin
				if(in == 0) begin
					state<=1028;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=4926;
					out<=17;
				end
				if(in == 3) begin
					state<=3008;
					out<=18;
				end
				if(in == 4) begin
					state<=6897;
					out<=19;
				end
			end
			1028: begin
				if(in == 0) begin
					state<=1029;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=4927;
					out<=22;
				end
				if(in == 3) begin
					state<=3009;
					out<=23;
				end
				if(in == 4) begin
					state<=6898;
					out<=24;
				end
			end
			1029: begin
				if(in == 0) begin
					state<=396;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=4294;
					out<=27;
				end
				if(in == 3) begin
					state<=3010;
					out<=28;
				end
				if(in == 4) begin
					state<=6899;
					out<=29;
				end
			end
			1030: begin
				if(in == 0) begin
					state<=1031;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=4929;
					out<=32;
				end
				if(in == 3) begin
					state<=3030;
					out<=33;
				end
				if(in == 4) begin
					state<=6919;
					out<=34;
				end
			end
			1031: begin
				if(in == 0) begin
					state<=1032;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=4930;
					out<=37;
				end
				if(in == 3) begin
					state<=3031;
					out<=38;
				end
				if(in == 4) begin
					state<=6920;
					out<=39;
				end
			end
			1032: begin
				if(in == 0) begin
					state<=1033;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=4931;
					out<=42;
				end
				if(in == 3) begin
					state<=3032;
					out<=43;
				end
				if(in == 4) begin
					state<=6921;
					out<=44;
				end
			end
			1033: begin
				if(in == 0) begin
					state<=1034;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=4932;
					out<=47;
				end
				if(in == 3) begin
					state<=3033;
					out<=48;
				end
				if(in == 4) begin
					state<=6922;
					out<=49;
				end
			end
			1034: begin
				if(in == 0) begin
					state<=1035;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=4933;
					out<=52;
				end
				if(in == 3) begin
					state<=3034;
					out<=53;
				end
				if(in == 4) begin
					state<=6923;
					out<=54;
				end
			end
			1035: begin
				if(in == 0) begin
					state<=1036;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=4934;
					out<=57;
				end
				if(in == 3) begin
					state<=3035;
					out<=58;
				end
				if(in == 4) begin
					state<=6924;
					out<=59;
				end
			end
			1036: begin
				if(in == 0) begin
					state<=1037;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=4935;
					out<=62;
				end
				if(in == 3) begin
					state<=3036;
					out<=63;
				end
				if(in == 4) begin
					state<=6925;
					out<=64;
				end
			end
			1037: begin
				if(in == 0) begin
					state<=1038;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=4936;
					out<=67;
				end
				if(in == 3) begin
					state<=3037;
					out<=68;
				end
				if(in == 4) begin
					state<=6926;
					out<=69;
				end
			end
			1038: begin
				if(in == 0) begin
					state<=1039;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=4937;
					out<=72;
				end
				if(in == 3) begin
					state<=3038;
					out<=73;
				end
				if(in == 4) begin
					state<=6927;
					out<=74;
				end
			end
			1039: begin
				if(in == 0) begin
					state<=1040;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=4938;
					out<=77;
				end
				if(in == 3) begin
					state<=3039;
					out<=78;
				end
				if(in == 4) begin
					state<=6928;
					out<=79;
				end
			end
			1040: begin
				if(in == 0) begin
					state<=1041;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=4939;
					out<=82;
				end
				if(in == 3) begin
					state<=3040;
					out<=83;
				end
				if(in == 4) begin
					state<=6929;
					out<=84;
				end
			end
			1041: begin
				if(in == 0) begin
					state<=1042;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=4940;
					out<=87;
				end
				if(in == 3) begin
					state<=3041;
					out<=88;
				end
				if(in == 4) begin
					state<=6930;
					out<=89;
				end
			end
			1042: begin
				if(in == 0) begin
					state<=1043;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=4941;
					out<=92;
				end
				if(in == 3) begin
					state<=3042;
					out<=93;
				end
				if(in == 4) begin
					state<=6931;
					out<=94;
				end
			end
			1043: begin
				if(in == 0) begin
					state<=1044;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=4942;
					out<=97;
				end
				if(in == 3) begin
					state<=3043;
					out<=98;
				end
				if(in == 4) begin
					state<=6932;
					out<=99;
				end
			end
			1044: begin
				if(in == 0) begin
					state<=1045;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=4943;
					out<=102;
				end
				if(in == 3) begin
					state<=3044;
					out<=103;
				end
				if(in == 4) begin
					state<=6933;
					out<=104;
				end
			end
			1045: begin
				if(in == 0) begin
					state<=1046;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=4944;
					out<=107;
				end
				if(in == 3) begin
					state<=3045;
					out<=108;
				end
				if(in == 4) begin
					state<=6934;
					out<=109;
				end
			end
			1046: begin
				if(in == 0) begin
					state<=1047;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=4945;
					out<=112;
				end
				if(in == 3) begin
					state<=3046;
					out<=113;
				end
				if(in == 4) begin
					state<=6935;
					out<=114;
				end
			end
			1047: begin
				if(in == 0) begin
					state<=1048;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=4946;
					out<=117;
				end
				if(in == 3) begin
					state<=3047;
					out<=118;
				end
				if(in == 4) begin
					state<=6936;
					out<=119;
				end
			end
			1048: begin
				if(in == 0) begin
					state<=1049;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=4947;
					out<=122;
				end
				if(in == 3) begin
					state<=3048;
					out<=123;
				end
				if(in == 4) begin
					state<=6937;
					out<=124;
				end
			end
			1049: begin
				if(in == 0) begin
					state<=1050;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=4948;
					out<=127;
				end
				if(in == 3) begin
					state<=3049;
					out<=128;
				end
				if(in == 4) begin
					state<=6938;
					out<=129;
				end
			end
			1050: begin
				if(in == 0) begin
					state<=1051;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=4949;
					out<=132;
				end
				if(in == 3) begin
					state<=3050;
					out<=133;
				end
				if(in == 4) begin
					state<=6939;
					out<=134;
				end
			end
			1051: begin
				if(in == 0) begin
					state<=1052;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=4950;
					out<=137;
				end
				if(in == 3) begin
					state<=3051;
					out<=138;
				end
				if(in == 4) begin
					state<=6940;
					out<=139;
				end
			end
			1052: begin
				if(in == 0) begin
					state<=1053;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=4951;
					out<=142;
				end
				if(in == 3) begin
					state<=3052;
					out<=143;
				end
				if(in == 4) begin
					state<=6941;
					out<=144;
				end
			end
			1053: begin
				if(in == 0) begin
					state<=1054;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=4952;
					out<=147;
				end
				if(in == 3) begin
					state<=3053;
					out<=148;
				end
				if(in == 4) begin
					state<=6942;
					out<=149;
				end
			end
			1054: begin
				if(in == 0) begin
					state<=1055;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=4953;
					out<=152;
				end
				if(in == 3) begin
					state<=3054;
					out<=153;
				end
				if(in == 4) begin
					state<=6943;
					out<=154;
				end
			end
			1055: begin
				if(in == 0) begin
					state<=1056;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=4954;
					out<=157;
				end
				if(in == 3) begin
					state<=3055;
					out<=158;
				end
				if(in == 4) begin
					state<=6944;
					out<=159;
				end
			end
			1056: begin
				if(in == 0) begin
					state<=1057;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=4955;
					out<=162;
				end
				if(in == 3) begin
					state<=3056;
					out<=163;
				end
				if(in == 4) begin
					state<=6945;
					out<=164;
				end
			end
			1057: begin
				if(in == 0) begin
					state<=1058;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=4956;
					out<=167;
				end
				if(in == 3) begin
					state<=3057;
					out<=168;
				end
				if(in == 4) begin
					state<=6946;
					out<=169;
				end
			end
			1058: begin
				if(in == 0) begin
					state<=1059;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=4957;
					out<=172;
				end
				if(in == 3) begin
					state<=3058;
					out<=173;
				end
				if(in == 4) begin
					state<=6947;
					out<=174;
				end
			end
			1059: begin
				if(in == 0) begin
					state<=1060;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=4958;
					out<=177;
				end
				if(in == 3) begin
					state<=3059;
					out<=178;
				end
				if(in == 4) begin
					state<=6948;
					out<=179;
				end
			end
			1060: begin
				if(in == 0) begin
					state<=1061;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=4959;
					out<=182;
				end
				if(in == 3) begin
					state<=3060;
					out<=183;
				end
				if(in == 4) begin
					state<=6949;
					out<=184;
				end
			end
			1061: begin
				if(in == 0) begin
					state<=1062;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=4960;
					out<=187;
				end
				if(in == 3) begin
					state<=3061;
					out<=188;
				end
				if(in == 4) begin
					state<=6950;
					out<=189;
				end
			end
			1062: begin
				if(in == 0) begin
					state<=1063;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=4961;
					out<=192;
				end
				if(in == 3) begin
					state<=3062;
					out<=193;
				end
				if(in == 4) begin
					state<=6951;
					out<=194;
				end
			end
			1063: begin
				if(in == 0) begin
					state<=1064;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=4962;
					out<=197;
				end
				if(in == 3) begin
					state<=3063;
					out<=198;
				end
				if(in == 4) begin
					state<=6952;
					out<=199;
				end
			end
			1064: begin
				if(in == 0) begin
					state<=1065;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=4963;
					out<=202;
				end
				if(in == 3) begin
					state<=3064;
					out<=203;
				end
				if(in == 4) begin
					state<=6953;
					out<=204;
				end
			end
			1065: begin
				if(in == 0) begin
					state<=1066;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=4964;
					out<=207;
				end
				if(in == 3) begin
					state<=3065;
					out<=208;
				end
				if(in == 4) begin
					state<=6954;
					out<=209;
				end
			end
			1066: begin
				if(in == 0) begin
					state<=1067;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=4965;
					out<=212;
				end
				if(in == 3) begin
					state<=3066;
					out<=213;
				end
				if(in == 4) begin
					state<=6955;
					out<=214;
				end
			end
			1067: begin
				if(in == 0) begin
					state<=1068;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=4966;
					out<=217;
				end
				if(in == 3) begin
					state<=3067;
					out<=218;
				end
				if(in == 4) begin
					state<=6956;
					out<=219;
				end
			end
			1068: begin
				if(in == 0) begin
					state<=1069;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=4967;
					out<=222;
				end
				if(in == 3) begin
					state<=3068;
					out<=223;
				end
				if(in == 4) begin
					state<=6957;
					out<=224;
				end
			end
			1069: begin
				if(in == 0) begin
					state<=1070;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=4968;
					out<=227;
				end
				if(in == 3) begin
					state<=3069;
					out<=228;
				end
				if(in == 4) begin
					state<=6958;
					out<=229;
				end
			end
			1070: begin
				if(in == 0) begin
					state<=1071;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=4969;
					out<=232;
				end
				if(in == 3) begin
					state<=3070;
					out<=233;
				end
				if(in == 4) begin
					state<=6959;
					out<=234;
				end
			end
			1071: begin
				if(in == 0) begin
					state<=1072;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=4970;
					out<=237;
				end
				if(in == 3) begin
					state<=3071;
					out<=238;
				end
				if(in == 4) begin
					state<=6960;
					out<=239;
				end
			end
			1072: begin
				if(in == 0) begin
					state<=1073;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=4971;
					out<=242;
				end
				if(in == 3) begin
					state<=3072;
					out<=243;
				end
				if(in == 4) begin
					state<=6961;
					out<=244;
				end
			end
			1073: begin
				if(in == 0) begin
					state<=1074;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=4972;
					out<=247;
				end
				if(in == 3) begin
					state<=3073;
					out<=248;
				end
				if(in == 4) begin
					state<=6962;
					out<=249;
				end
			end
			1074: begin
				if(in == 0) begin
					state<=1075;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=4973;
					out<=252;
				end
				if(in == 3) begin
					state<=3074;
					out<=253;
				end
				if(in == 4) begin
					state<=6963;
					out<=254;
				end
			end
			1075: begin
				if(in == 0) begin
					state<=1076;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=4974;
					out<=1;
				end
				if(in == 3) begin
					state<=3075;
					out<=2;
				end
				if(in == 4) begin
					state<=6964;
					out<=3;
				end
			end
			1076: begin
				if(in == 0) begin
					state<=1077;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=4975;
					out<=6;
				end
				if(in == 3) begin
					state<=3076;
					out<=7;
				end
				if(in == 4) begin
					state<=6965;
					out<=8;
				end
			end
			1077: begin
				if(in == 0) begin
					state<=1078;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=4976;
					out<=11;
				end
				if(in == 3) begin
					state<=3077;
					out<=12;
				end
				if(in == 4) begin
					state<=6966;
					out<=13;
				end
			end
			1078: begin
				if(in == 0) begin
					state<=1079;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=4977;
					out<=16;
				end
				if(in == 3) begin
					state<=3078;
					out<=17;
				end
				if(in == 4) begin
					state<=6967;
					out<=18;
				end
			end
			1079: begin
				if(in == 0) begin
					state<=1080;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=4978;
					out<=21;
				end
				if(in == 3) begin
					state<=3079;
					out<=22;
				end
				if(in == 4) begin
					state<=6968;
					out<=23;
				end
			end
			1080: begin
				if(in == 0) begin
					state<=1081;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=4979;
					out<=26;
				end
				if(in == 3) begin
					state<=3080;
					out<=27;
				end
				if(in == 4) begin
					state<=6969;
					out<=28;
				end
			end
			1081: begin
				if(in == 0) begin
					state<=1082;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=4980;
					out<=31;
				end
				if(in == 3) begin
					state<=3081;
					out<=32;
				end
				if(in == 4) begin
					state<=6970;
					out<=33;
				end
			end
			1082: begin
				if(in == 0) begin
					state<=1083;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=4981;
					out<=36;
				end
				if(in == 3) begin
					state<=3082;
					out<=37;
				end
				if(in == 4) begin
					state<=6971;
					out<=38;
				end
			end
			1083: begin
				if(in == 0) begin
					state<=1084;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=4982;
					out<=41;
				end
				if(in == 3) begin
					state<=3083;
					out<=42;
				end
				if(in == 4) begin
					state<=6972;
					out<=43;
				end
			end
			1084: begin
				if(in == 0) begin
					state<=1085;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=4983;
					out<=46;
				end
				if(in == 3) begin
					state<=3084;
					out<=47;
				end
				if(in == 4) begin
					state<=6973;
					out<=48;
				end
			end
			1085: begin
				if(in == 0) begin
					state<=1086;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=4984;
					out<=51;
				end
				if(in == 3) begin
					state<=3085;
					out<=52;
				end
				if(in == 4) begin
					state<=6974;
					out<=53;
				end
			end
			1086: begin
				if(in == 0) begin
					state<=1087;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=4985;
					out<=56;
				end
				if(in == 3) begin
					state<=3086;
					out<=57;
				end
				if(in == 4) begin
					state<=6975;
					out<=58;
				end
			end
			1087: begin
				if(in == 0) begin
					state<=1088;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=4986;
					out<=61;
				end
				if(in == 3) begin
					state<=3087;
					out<=62;
				end
				if(in == 4) begin
					state<=6976;
					out<=63;
				end
			end
			1088: begin
				if(in == 0) begin
					state<=1089;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=4987;
					out<=66;
				end
				if(in == 3) begin
					state<=3088;
					out<=67;
				end
				if(in == 4) begin
					state<=6977;
					out<=68;
				end
			end
			1089: begin
				if(in == 0) begin
					state<=1090;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=4988;
					out<=71;
				end
				if(in == 3) begin
					state<=3089;
					out<=72;
				end
				if(in == 4) begin
					state<=6978;
					out<=73;
				end
			end
			1090: begin
				if(in == 0) begin
					state<=1091;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=4989;
					out<=76;
				end
				if(in == 3) begin
					state<=3090;
					out<=77;
				end
				if(in == 4) begin
					state<=6979;
					out<=78;
				end
			end
			1091: begin
				if(in == 0) begin
					state<=1092;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=4990;
					out<=81;
				end
				if(in == 3) begin
					state<=3091;
					out<=82;
				end
				if(in == 4) begin
					state<=6980;
					out<=83;
				end
			end
			1092: begin
				if(in == 0) begin
					state<=1093;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=4991;
					out<=86;
				end
				if(in == 3) begin
					state<=3092;
					out<=87;
				end
				if(in == 4) begin
					state<=6981;
					out<=88;
				end
			end
			1093: begin
				if(in == 0) begin
					state<=1094;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=4992;
					out<=91;
				end
				if(in == 3) begin
					state<=3093;
					out<=92;
				end
				if(in == 4) begin
					state<=6982;
					out<=93;
				end
			end
			1094: begin
				if(in == 0) begin
					state<=1095;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=4993;
					out<=96;
				end
				if(in == 3) begin
					state<=3094;
					out<=97;
				end
				if(in == 4) begin
					state<=6983;
					out<=98;
				end
			end
			1095: begin
				if(in == 0) begin
					state<=1096;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=4994;
					out<=101;
				end
				if(in == 3) begin
					state<=3095;
					out<=102;
				end
				if(in == 4) begin
					state<=6984;
					out<=103;
				end
			end
			1096: begin
				if(in == 0) begin
					state<=1097;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=4995;
					out<=106;
				end
				if(in == 3) begin
					state<=3096;
					out<=107;
				end
				if(in == 4) begin
					state<=6985;
					out<=108;
				end
			end
			1097: begin
				if(in == 0) begin
					state<=1098;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=4996;
					out<=111;
				end
				if(in == 3) begin
					state<=3097;
					out<=112;
				end
				if(in == 4) begin
					state<=6986;
					out<=113;
				end
			end
			1098: begin
				if(in == 0) begin
					state<=1099;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=4997;
					out<=116;
				end
				if(in == 3) begin
					state<=3098;
					out<=117;
				end
				if(in == 4) begin
					state<=6987;
					out<=118;
				end
			end
			1099: begin
				if(in == 0) begin
					state<=1100;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=4998;
					out<=121;
				end
				if(in == 3) begin
					state<=3099;
					out<=122;
				end
				if(in == 4) begin
					state<=6988;
					out<=123;
				end
			end
			1100: begin
				if(in == 0) begin
					state<=1101;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=4999;
					out<=126;
				end
				if(in == 3) begin
					state<=3100;
					out<=127;
				end
				if(in == 4) begin
					state<=6989;
					out<=128;
				end
			end
			1101: begin
				if(in == 0) begin
					state<=1102;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=5000;
					out<=131;
				end
				if(in == 3) begin
					state<=3101;
					out<=132;
				end
				if(in == 4) begin
					state<=6990;
					out<=133;
				end
			end
			1102: begin
				if(in == 0) begin
					state<=1103;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=5001;
					out<=136;
				end
				if(in == 3) begin
					state<=3102;
					out<=137;
				end
				if(in == 4) begin
					state<=6991;
					out<=138;
				end
			end
			1103: begin
				if(in == 0) begin
					state<=1104;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=5002;
					out<=141;
				end
				if(in == 3) begin
					state<=3103;
					out<=142;
				end
				if(in == 4) begin
					state<=6992;
					out<=143;
				end
			end
			1104: begin
				if(in == 0) begin
					state<=1105;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=5003;
					out<=146;
				end
				if(in == 3) begin
					state<=3104;
					out<=147;
				end
				if(in == 4) begin
					state<=6993;
					out<=148;
				end
			end
			1105: begin
				if(in == 0) begin
					state<=1106;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=5004;
					out<=151;
				end
				if(in == 3) begin
					state<=3105;
					out<=152;
				end
				if(in == 4) begin
					state<=6994;
					out<=153;
				end
			end
			1106: begin
				if(in == 0) begin
					state<=1107;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=5005;
					out<=156;
				end
				if(in == 3) begin
					state<=3106;
					out<=157;
				end
				if(in == 4) begin
					state<=6995;
					out<=158;
				end
			end
			1107: begin
				if(in == 0) begin
					state<=1108;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=5006;
					out<=161;
				end
				if(in == 3) begin
					state<=3107;
					out<=162;
				end
				if(in == 4) begin
					state<=6996;
					out<=163;
				end
			end
			1108: begin
				if(in == 0) begin
					state<=1109;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=5007;
					out<=166;
				end
				if(in == 3) begin
					state<=3108;
					out<=167;
				end
				if(in == 4) begin
					state<=6997;
					out<=168;
				end
			end
			1109: begin
				if(in == 0) begin
					state<=1110;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=5008;
					out<=171;
				end
				if(in == 3) begin
					state<=3109;
					out<=172;
				end
				if(in == 4) begin
					state<=6998;
					out<=173;
				end
			end
			1110: begin
				if(in == 0) begin
					state<=1111;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=5009;
					out<=176;
				end
				if(in == 3) begin
					state<=3110;
					out<=177;
				end
				if(in == 4) begin
					state<=6999;
					out<=178;
				end
			end
			1111: begin
				if(in == 0) begin
					state<=1112;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=5010;
					out<=181;
				end
				if(in == 3) begin
					state<=3111;
					out<=182;
				end
				if(in == 4) begin
					state<=7000;
					out<=183;
				end
			end
			1112: begin
				if(in == 0) begin
					state<=1113;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=5011;
					out<=186;
				end
				if(in == 3) begin
					state<=3112;
					out<=187;
				end
				if(in == 4) begin
					state<=7001;
					out<=188;
				end
			end
			1113: begin
				if(in == 0) begin
					state<=1114;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=5012;
					out<=191;
				end
				if(in == 3) begin
					state<=3113;
					out<=192;
				end
				if(in == 4) begin
					state<=7002;
					out<=193;
				end
			end
			1114: begin
				if(in == 0) begin
					state<=1115;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=5013;
					out<=196;
				end
				if(in == 3) begin
					state<=3114;
					out<=197;
				end
				if(in == 4) begin
					state<=7003;
					out<=198;
				end
			end
			1115: begin
				if(in == 0) begin
					state<=1116;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=5014;
					out<=201;
				end
				if(in == 3) begin
					state<=3115;
					out<=202;
				end
				if(in == 4) begin
					state<=7004;
					out<=203;
				end
			end
			1116: begin
				if(in == 0) begin
					state<=1117;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=5015;
					out<=206;
				end
				if(in == 3) begin
					state<=3116;
					out<=207;
				end
				if(in == 4) begin
					state<=7005;
					out<=208;
				end
			end
			1117: begin
				if(in == 0) begin
					state<=1118;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=5016;
					out<=211;
				end
				if(in == 3) begin
					state<=3117;
					out<=212;
				end
				if(in == 4) begin
					state<=7006;
					out<=213;
				end
			end
			1118: begin
				if(in == 0) begin
					state<=1119;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=5017;
					out<=216;
				end
				if(in == 3) begin
					state<=3118;
					out<=217;
				end
				if(in == 4) begin
					state<=7007;
					out<=218;
				end
			end
			1119: begin
				if(in == 0) begin
					state<=1120;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=5018;
					out<=221;
				end
				if(in == 3) begin
					state<=3119;
					out<=222;
				end
				if(in == 4) begin
					state<=7008;
					out<=223;
				end
			end
			1120: begin
				if(in == 0) begin
					state<=1121;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=5019;
					out<=226;
				end
				if(in == 3) begin
					state<=3120;
					out<=227;
				end
				if(in == 4) begin
					state<=7009;
					out<=228;
				end
			end
			1121: begin
				if(in == 0) begin
					state<=1122;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=5020;
					out<=231;
				end
				if(in == 3) begin
					state<=3121;
					out<=232;
				end
				if(in == 4) begin
					state<=7010;
					out<=233;
				end
			end
			1122: begin
				if(in == 0) begin
					state<=1123;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=5021;
					out<=236;
				end
				if(in == 3) begin
					state<=3122;
					out<=237;
				end
				if(in == 4) begin
					state<=7011;
					out<=238;
				end
			end
			1123: begin
				if(in == 0) begin
					state<=1124;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=5022;
					out<=241;
				end
				if(in == 3) begin
					state<=3123;
					out<=242;
				end
				if(in == 4) begin
					state<=7012;
					out<=243;
				end
			end
			1124: begin
				if(in == 0) begin
					state<=1125;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=5023;
					out<=246;
				end
				if(in == 3) begin
					state<=3124;
					out<=247;
				end
				if(in == 4) begin
					state<=7013;
					out<=248;
				end
			end
			1125: begin
				if(in == 0) begin
					state<=1126;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=5024;
					out<=251;
				end
				if(in == 3) begin
					state<=3125;
					out<=252;
				end
				if(in == 4) begin
					state<=7014;
					out<=253;
				end
			end
			1126: begin
				if(in == 0) begin
					state<=1127;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=5025;
					out<=0;
				end
				if(in == 3) begin
					state<=3126;
					out<=1;
				end
				if(in == 4) begin
					state<=7015;
					out<=2;
				end
			end
			1127: begin
				if(in == 0) begin
					state<=1128;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=5026;
					out<=5;
				end
				if(in == 3) begin
					state<=3127;
					out<=6;
				end
				if(in == 4) begin
					state<=7016;
					out<=7;
				end
			end
			1128: begin
				if(in == 0) begin
					state<=1129;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=5027;
					out<=10;
				end
				if(in == 3) begin
					state<=3128;
					out<=11;
				end
				if(in == 4) begin
					state<=7017;
					out<=12;
				end
			end
			1129: begin
				if(in == 0) begin
					state<=1130;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=5028;
					out<=15;
				end
				if(in == 3) begin
					state<=3129;
					out<=16;
				end
				if(in == 4) begin
					state<=7018;
					out<=17;
				end
			end
			1130: begin
				if(in == 0) begin
					state<=1131;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=5029;
					out<=20;
				end
				if(in == 3) begin
					state<=3130;
					out<=21;
				end
				if(in == 4) begin
					state<=7019;
					out<=22;
				end
			end
			1131: begin
				if(in == 0) begin
					state<=1132;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=5030;
					out<=25;
				end
				if(in == 3) begin
					state<=3131;
					out<=26;
				end
				if(in == 4) begin
					state<=7020;
					out<=27;
				end
			end
			1132: begin
				if(in == 0) begin
					state<=1133;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=5031;
					out<=30;
				end
				if(in == 3) begin
					state<=3132;
					out<=31;
				end
				if(in == 4) begin
					state<=7021;
					out<=32;
				end
			end
			1133: begin
				if(in == 0) begin
					state<=1134;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=5032;
					out<=35;
				end
				if(in == 3) begin
					state<=3133;
					out<=36;
				end
				if(in == 4) begin
					state<=7022;
					out<=37;
				end
			end
			1134: begin
				if(in == 0) begin
					state<=1135;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=5033;
					out<=40;
				end
				if(in == 3) begin
					state<=3134;
					out<=41;
				end
				if(in == 4) begin
					state<=7023;
					out<=42;
				end
			end
			1135: begin
				if(in == 0) begin
					state<=1136;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=5034;
					out<=45;
				end
				if(in == 3) begin
					state<=3135;
					out<=46;
				end
				if(in == 4) begin
					state<=7024;
					out<=47;
				end
			end
			1136: begin
				if(in == 0) begin
					state<=1137;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=5035;
					out<=50;
				end
				if(in == 3) begin
					state<=3136;
					out<=51;
				end
				if(in == 4) begin
					state<=7025;
					out<=52;
				end
			end
			1137: begin
				if(in == 0) begin
					state<=1138;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=5036;
					out<=55;
				end
				if(in == 3) begin
					state<=3137;
					out<=56;
				end
				if(in == 4) begin
					state<=7026;
					out<=57;
				end
			end
			1138: begin
				if(in == 0) begin
					state<=1139;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=5037;
					out<=60;
				end
				if(in == 3) begin
					state<=3138;
					out<=61;
				end
				if(in == 4) begin
					state<=7027;
					out<=62;
				end
			end
			1139: begin
				if(in == 0) begin
					state<=1140;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=5038;
					out<=65;
				end
				if(in == 3) begin
					state<=3139;
					out<=66;
				end
				if(in == 4) begin
					state<=7028;
					out<=67;
				end
			end
			1140: begin
				if(in == 0) begin
					state<=1141;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=5039;
					out<=70;
				end
				if(in == 3) begin
					state<=3140;
					out<=71;
				end
				if(in == 4) begin
					state<=7029;
					out<=72;
				end
			end
			1141: begin
				if(in == 0) begin
					state<=1142;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=5040;
					out<=75;
				end
				if(in == 3) begin
					state<=3141;
					out<=76;
				end
				if(in == 4) begin
					state<=7030;
					out<=77;
				end
			end
			1142: begin
				if(in == 0) begin
					state<=1143;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=5041;
					out<=80;
				end
				if(in == 3) begin
					state<=3142;
					out<=81;
				end
				if(in == 4) begin
					state<=7031;
					out<=82;
				end
			end
			1143: begin
				if(in == 0) begin
					state<=1144;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=5042;
					out<=85;
				end
				if(in == 3) begin
					state<=3143;
					out<=86;
				end
				if(in == 4) begin
					state<=7032;
					out<=87;
				end
			end
			1144: begin
				if(in == 0) begin
					state<=1145;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=5043;
					out<=90;
				end
				if(in == 3) begin
					state<=3144;
					out<=91;
				end
				if(in == 4) begin
					state<=7033;
					out<=92;
				end
			end
			1145: begin
				if(in == 0) begin
					state<=1146;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=5044;
					out<=95;
				end
				if(in == 3) begin
					state<=3145;
					out<=96;
				end
				if(in == 4) begin
					state<=7034;
					out<=97;
				end
			end
			1146: begin
				if(in == 0) begin
					state<=1147;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=5045;
					out<=100;
				end
				if(in == 3) begin
					state<=3146;
					out<=101;
				end
				if(in == 4) begin
					state<=7035;
					out<=102;
				end
			end
			1147: begin
				if(in == 0) begin
					state<=1148;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=5046;
					out<=105;
				end
				if(in == 3) begin
					state<=3147;
					out<=106;
				end
				if(in == 4) begin
					state<=7036;
					out<=107;
				end
			end
			1148: begin
				if(in == 0) begin
					state<=1149;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=5047;
					out<=110;
				end
				if(in == 3) begin
					state<=3148;
					out<=111;
				end
				if(in == 4) begin
					state<=7037;
					out<=112;
				end
			end
			1149: begin
				if(in == 0) begin
					state<=1150;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=5048;
					out<=115;
				end
				if(in == 3) begin
					state<=3149;
					out<=116;
				end
				if(in == 4) begin
					state<=7038;
					out<=117;
				end
			end
			1150: begin
				if(in == 0) begin
					state<=1151;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=5049;
					out<=120;
				end
				if(in == 3) begin
					state<=3150;
					out<=121;
				end
				if(in == 4) begin
					state<=7039;
					out<=122;
				end
			end
			1151: begin
				if(in == 0) begin
					state<=1152;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=5050;
					out<=125;
				end
				if(in == 3) begin
					state<=3151;
					out<=126;
				end
				if(in == 4) begin
					state<=7040;
					out<=127;
				end
			end
			1152: begin
				if(in == 0) begin
					state<=1153;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=5051;
					out<=130;
				end
				if(in == 3) begin
					state<=3152;
					out<=131;
				end
				if(in == 4) begin
					state<=7041;
					out<=132;
				end
			end
			1153: begin
				if(in == 0) begin
					state<=1154;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=5052;
					out<=135;
				end
				if(in == 3) begin
					state<=3153;
					out<=136;
				end
				if(in == 4) begin
					state<=7042;
					out<=137;
				end
			end
			1154: begin
				if(in == 0) begin
					state<=1155;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=5053;
					out<=140;
				end
				if(in == 3) begin
					state<=3154;
					out<=141;
				end
				if(in == 4) begin
					state<=7043;
					out<=142;
				end
			end
			1155: begin
				if(in == 0) begin
					state<=1156;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=5054;
					out<=145;
				end
				if(in == 3) begin
					state<=3155;
					out<=146;
				end
				if(in == 4) begin
					state<=7044;
					out<=147;
				end
			end
			1156: begin
				if(in == 0) begin
					state<=1157;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=5055;
					out<=150;
				end
				if(in == 3) begin
					state<=3156;
					out<=151;
				end
				if(in == 4) begin
					state<=7045;
					out<=152;
				end
			end
			1157: begin
				if(in == 0) begin
					state<=1158;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=5056;
					out<=155;
				end
				if(in == 3) begin
					state<=3157;
					out<=156;
				end
				if(in == 4) begin
					state<=7046;
					out<=157;
				end
			end
			1158: begin
				if(in == 0) begin
					state<=1159;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=5057;
					out<=160;
				end
				if(in == 3) begin
					state<=3158;
					out<=161;
				end
				if(in == 4) begin
					state<=7047;
					out<=162;
				end
			end
			1159: begin
				if(in == 0) begin
					state<=1160;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=5058;
					out<=165;
				end
				if(in == 3) begin
					state<=3159;
					out<=166;
				end
				if(in == 4) begin
					state<=7048;
					out<=167;
				end
			end
			1160: begin
				if(in == 0) begin
					state<=1161;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=5059;
					out<=170;
				end
				if(in == 3) begin
					state<=3160;
					out<=171;
				end
				if(in == 4) begin
					state<=7049;
					out<=172;
				end
			end
			1161: begin
				if(in == 0) begin
					state<=1162;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=5060;
					out<=175;
				end
				if(in == 3) begin
					state<=3161;
					out<=176;
				end
				if(in == 4) begin
					state<=7050;
					out<=177;
				end
			end
			1162: begin
				if(in == 0) begin
					state<=1163;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=5061;
					out<=180;
				end
				if(in == 3) begin
					state<=3162;
					out<=181;
				end
				if(in == 4) begin
					state<=7051;
					out<=182;
				end
			end
			1163: begin
				if(in == 0) begin
					state<=1164;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=5062;
					out<=185;
				end
				if(in == 3) begin
					state<=3163;
					out<=186;
				end
				if(in == 4) begin
					state<=7052;
					out<=187;
				end
			end
			1164: begin
				if(in == 0) begin
					state<=1165;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=5063;
					out<=190;
				end
				if(in == 3) begin
					state<=3164;
					out<=191;
				end
				if(in == 4) begin
					state<=7053;
					out<=192;
				end
			end
			1165: begin
				if(in == 0) begin
					state<=1166;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=5064;
					out<=195;
				end
				if(in == 3) begin
					state<=3165;
					out<=196;
				end
				if(in == 4) begin
					state<=7054;
					out<=197;
				end
			end
			1166: begin
				if(in == 0) begin
					state<=1167;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=5065;
					out<=200;
				end
				if(in == 3) begin
					state<=3166;
					out<=201;
				end
				if(in == 4) begin
					state<=7055;
					out<=202;
				end
			end
			1167: begin
				if(in == 0) begin
					state<=1168;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=5066;
					out<=205;
				end
				if(in == 3) begin
					state<=3167;
					out<=206;
				end
				if(in == 4) begin
					state<=7056;
					out<=207;
				end
			end
			1168: begin
				if(in == 0) begin
					state<=1169;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=5067;
					out<=210;
				end
				if(in == 3) begin
					state<=3168;
					out<=211;
				end
				if(in == 4) begin
					state<=7057;
					out<=212;
				end
			end
			1169: begin
				if(in == 0) begin
					state<=1170;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=5068;
					out<=215;
				end
				if(in == 3) begin
					state<=3169;
					out<=216;
				end
				if(in == 4) begin
					state<=7058;
					out<=217;
				end
			end
			1170: begin
				if(in == 0) begin
					state<=1171;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=5069;
					out<=220;
				end
				if(in == 3) begin
					state<=3170;
					out<=221;
				end
				if(in == 4) begin
					state<=7059;
					out<=222;
				end
			end
			1171: begin
				if(in == 0) begin
					state<=1172;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=5070;
					out<=225;
				end
				if(in == 3) begin
					state<=3171;
					out<=226;
				end
				if(in == 4) begin
					state<=7060;
					out<=227;
				end
			end
			1172: begin
				if(in == 0) begin
					state<=1173;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=5071;
					out<=230;
				end
				if(in == 3) begin
					state<=3172;
					out<=231;
				end
				if(in == 4) begin
					state<=7061;
					out<=232;
				end
			end
			1173: begin
				if(in == 0) begin
					state<=1174;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=5072;
					out<=235;
				end
				if(in == 3) begin
					state<=3173;
					out<=236;
				end
				if(in == 4) begin
					state<=7062;
					out<=237;
				end
			end
			1174: begin
				if(in == 0) begin
					state<=1175;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=5073;
					out<=240;
				end
				if(in == 3) begin
					state<=3174;
					out<=241;
				end
				if(in == 4) begin
					state<=7063;
					out<=242;
				end
			end
			1175: begin
				if(in == 0) begin
					state<=1176;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=5074;
					out<=245;
				end
				if(in == 3) begin
					state<=3175;
					out<=246;
				end
				if(in == 4) begin
					state<=7064;
					out<=247;
				end
			end
			1176: begin
				if(in == 0) begin
					state<=1177;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=5075;
					out<=250;
				end
				if(in == 3) begin
					state<=3176;
					out<=251;
				end
				if(in == 4) begin
					state<=7065;
					out<=252;
				end
			end
			1177: begin
				if(in == 0) begin
					state<=1178;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=5076;
					out<=255;
				end
				if(in == 3) begin
					state<=3177;
					out<=0;
				end
				if(in == 4) begin
					state<=7066;
					out<=1;
				end
			end
			1178: begin
				if(in == 0) begin
					state<=1179;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=5077;
					out<=4;
				end
				if(in == 3) begin
					state<=3178;
					out<=5;
				end
				if(in == 4) begin
					state<=7067;
					out<=6;
				end
			end
			1179: begin
				if(in == 0) begin
					state<=1180;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=5078;
					out<=9;
				end
				if(in == 3) begin
					state<=3179;
					out<=10;
				end
				if(in == 4) begin
					state<=7068;
					out<=11;
				end
			end
			1180: begin
				if(in == 0) begin
					state<=1181;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=5079;
					out<=14;
				end
				if(in == 3) begin
					state<=3180;
					out<=15;
				end
				if(in == 4) begin
					state<=7069;
					out<=16;
				end
			end
			1181: begin
				if(in == 0) begin
					state<=1182;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=5080;
					out<=19;
				end
				if(in == 3) begin
					state<=3181;
					out<=20;
				end
				if(in == 4) begin
					state<=7070;
					out<=21;
				end
			end
			1182: begin
				if(in == 0) begin
					state<=1183;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=5081;
					out<=24;
				end
				if(in == 3) begin
					state<=3182;
					out<=25;
				end
				if(in == 4) begin
					state<=7071;
					out<=26;
				end
			end
			1183: begin
				if(in == 0) begin
					state<=1184;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=5082;
					out<=29;
				end
				if(in == 3) begin
					state<=3183;
					out<=30;
				end
				if(in == 4) begin
					state<=7072;
					out<=31;
				end
			end
			1184: begin
				if(in == 0) begin
					state<=1185;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=5083;
					out<=34;
				end
				if(in == 3) begin
					state<=3184;
					out<=35;
				end
				if(in == 4) begin
					state<=7073;
					out<=36;
				end
			end
			1185: begin
				if(in == 0) begin
					state<=1186;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=5084;
					out<=39;
				end
				if(in == 3) begin
					state<=3185;
					out<=40;
				end
				if(in == 4) begin
					state<=7074;
					out<=41;
				end
			end
			1186: begin
				if(in == 0) begin
					state<=1187;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=5085;
					out<=44;
				end
				if(in == 3) begin
					state<=3186;
					out<=45;
				end
				if(in == 4) begin
					state<=7075;
					out<=46;
				end
			end
			1187: begin
				if(in == 0) begin
					state<=1188;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=5086;
					out<=49;
				end
				if(in == 3) begin
					state<=3187;
					out<=50;
				end
				if(in == 4) begin
					state<=7076;
					out<=51;
				end
			end
			1188: begin
				if(in == 0) begin
					state<=1189;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=5087;
					out<=54;
				end
				if(in == 3) begin
					state<=3188;
					out<=55;
				end
				if(in == 4) begin
					state<=7077;
					out<=56;
				end
			end
			1189: begin
				if(in == 0) begin
					state<=1190;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=5088;
					out<=59;
				end
				if(in == 3) begin
					state<=3189;
					out<=60;
				end
				if(in == 4) begin
					state<=7078;
					out<=61;
				end
			end
			1190: begin
				if(in == 0) begin
					state<=1191;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=5089;
					out<=64;
				end
				if(in == 3) begin
					state<=3190;
					out<=65;
				end
				if(in == 4) begin
					state<=7079;
					out<=66;
				end
			end
			1191: begin
				if(in == 0) begin
					state<=1192;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=5090;
					out<=69;
				end
				if(in == 3) begin
					state<=3191;
					out<=70;
				end
				if(in == 4) begin
					state<=7080;
					out<=71;
				end
			end
			1192: begin
				if(in == 0) begin
					state<=1193;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=5091;
					out<=74;
				end
				if(in == 3) begin
					state<=3192;
					out<=75;
				end
				if(in == 4) begin
					state<=7081;
					out<=76;
				end
			end
			1193: begin
				if(in == 0) begin
					state<=1194;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=5092;
					out<=79;
				end
				if(in == 3) begin
					state<=3193;
					out<=80;
				end
				if(in == 4) begin
					state<=7082;
					out<=81;
				end
			end
			1194: begin
				if(in == 0) begin
					state<=1195;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=5093;
					out<=84;
				end
				if(in == 3) begin
					state<=3194;
					out<=85;
				end
				if(in == 4) begin
					state<=7083;
					out<=86;
				end
			end
			1195: begin
				if(in == 0) begin
					state<=1196;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=5094;
					out<=89;
				end
				if(in == 3) begin
					state<=3195;
					out<=90;
				end
				if(in == 4) begin
					state<=7084;
					out<=91;
				end
			end
			1196: begin
				if(in == 0) begin
					state<=1197;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=5095;
					out<=94;
				end
				if(in == 3) begin
					state<=3196;
					out<=95;
				end
				if(in == 4) begin
					state<=7085;
					out<=96;
				end
			end
			1197: begin
				if(in == 0) begin
					state<=1198;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=5096;
					out<=99;
				end
				if(in == 3) begin
					state<=3197;
					out<=100;
				end
				if(in == 4) begin
					state<=7086;
					out<=101;
				end
			end
			1198: begin
				if(in == 0) begin
					state<=1199;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=5097;
					out<=104;
				end
				if(in == 3) begin
					state<=3198;
					out<=105;
				end
				if(in == 4) begin
					state<=7087;
					out<=106;
				end
			end
			1199: begin
				if(in == 0) begin
					state<=1200;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=5098;
					out<=109;
				end
				if(in == 3) begin
					state<=3199;
					out<=110;
				end
				if(in == 4) begin
					state<=7088;
					out<=111;
				end
			end
			1200: begin
				if(in == 0) begin
					state<=1201;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=5099;
					out<=114;
				end
				if(in == 3) begin
					state<=3200;
					out<=115;
				end
				if(in == 4) begin
					state<=7089;
					out<=116;
				end
			end
			1201: begin
				if(in == 0) begin
					state<=1202;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=5100;
					out<=119;
				end
				if(in == 3) begin
					state<=3201;
					out<=120;
				end
				if(in == 4) begin
					state<=7090;
					out<=121;
				end
			end
			1202: begin
				if(in == 0) begin
					state<=1203;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=5101;
					out<=124;
				end
				if(in == 3) begin
					state<=3202;
					out<=125;
				end
				if(in == 4) begin
					state<=7091;
					out<=126;
				end
			end
			1203: begin
				if(in == 0) begin
					state<=1204;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=5102;
					out<=129;
				end
				if(in == 3) begin
					state<=3203;
					out<=130;
				end
				if(in == 4) begin
					state<=7092;
					out<=131;
				end
			end
			1204: begin
				if(in == 0) begin
					state<=1205;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=5103;
					out<=134;
				end
				if(in == 3) begin
					state<=3204;
					out<=135;
				end
				if(in == 4) begin
					state<=7093;
					out<=136;
				end
			end
			1205: begin
				if(in == 0) begin
					state<=1206;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=5104;
					out<=139;
				end
				if(in == 3) begin
					state<=3205;
					out<=140;
				end
				if(in == 4) begin
					state<=7094;
					out<=141;
				end
			end
			1206: begin
				if(in == 0) begin
					state<=1207;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=5105;
					out<=144;
				end
				if(in == 3) begin
					state<=3206;
					out<=145;
				end
				if(in == 4) begin
					state<=7095;
					out<=146;
				end
			end
			1207: begin
				if(in == 0) begin
					state<=1208;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=5106;
					out<=149;
				end
				if(in == 3) begin
					state<=3207;
					out<=150;
				end
				if(in == 4) begin
					state<=7096;
					out<=151;
				end
			end
			1208: begin
				if(in == 0) begin
					state<=1209;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=5107;
					out<=154;
				end
				if(in == 3) begin
					state<=3208;
					out<=155;
				end
				if(in == 4) begin
					state<=7097;
					out<=156;
				end
			end
			1209: begin
				if(in == 0) begin
					state<=1210;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=5108;
					out<=159;
				end
				if(in == 3) begin
					state<=3209;
					out<=160;
				end
				if(in == 4) begin
					state<=7098;
					out<=161;
				end
			end
			1210: begin
				if(in == 0) begin
					state<=1211;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=5109;
					out<=164;
				end
				if(in == 3) begin
					state<=3210;
					out<=165;
				end
				if(in == 4) begin
					state<=7099;
					out<=166;
				end
			end
			1211: begin
				if(in == 0) begin
					state<=1212;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=5110;
					out<=169;
				end
				if(in == 3) begin
					state<=3211;
					out<=170;
				end
				if(in == 4) begin
					state<=7100;
					out<=171;
				end
			end
			1212: begin
				if(in == 0) begin
					state<=1213;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=5111;
					out<=174;
				end
				if(in == 3) begin
					state<=3212;
					out<=175;
				end
				if(in == 4) begin
					state<=7101;
					out<=176;
				end
			end
			1213: begin
				if(in == 0) begin
					state<=1214;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=5112;
					out<=179;
				end
				if(in == 3) begin
					state<=3213;
					out<=180;
				end
				if(in == 4) begin
					state<=7102;
					out<=181;
				end
			end
			1214: begin
				if(in == 0) begin
					state<=1215;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=5113;
					out<=184;
				end
				if(in == 3) begin
					state<=3214;
					out<=185;
				end
				if(in == 4) begin
					state<=7103;
					out<=186;
				end
			end
			1215: begin
				if(in == 0) begin
					state<=1216;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=5114;
					out<=189;
				end
				if(in == 3) begin
					state<=3215;
					out<=190;
				end
				if(in == 4) begin
					state<=7104;
					out<=191;
				end
			end
			1216: begin
				if(in == 0) begin
					state<=1217;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=5115;
					out<=194;
				end
				if(in == 3) begin
					state<=3216;
					out<=195;
				end
				if(in == 4) begin
					state<=7105;
					out<=196;
				end
			end
			1217: begin
				if(in == 0) begin
					state<=1218;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=5116;
					out<=199;
				end
				if(in == 3) begin
					state<=3217;
					out<=200;
				end
				if(in == 4) begin
					state<=7106;
					out<=201;
				end
			end
			1218: begin
				if(in == 0) begin
					state<=1219;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=5117;
					out<=204;
				end
				if(in == 3) begin
					state<=3218;
					out<=205;
				end
				if(in == 4) begin
					state<=7107;
					out<=206;
				end
			end
			1219: begin
				if(in == 0) begin
					state<=1220;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=5118;
					out<=209;
				end
				if(in == 3) begin
					state<=3219;
					out<=210;
				end
				if(in == 4) begin
					state<=7108;
					out<=211;
				end
			end
			1220: begin
				if(in == 0) begin
					state<=1221;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=5119;
					out<=214;
				end
				if(in == 3) begin
					state<=3220;
					out<=215;
				end
				if(in == 4) begin
					state<=7109;
					out<=216;
				end
			end
			1221: begin
				if(in == 0) begin
					state<=1222;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=5120;
					out<=219;
				end
				if(in == 3) begin
					state<=3221;
					out<=220;
				end
				if(in == 4) begin
					state<=7110;
					out<=221;
				end
			end
			1222: begin
				if(in == 0) begin
					state<=1223;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=5121;
					out<=224;
				end
				if(in == 3) begin
					state<=3222;
					out<=225;
				end
				if(in == 4) begin
					state<=7111;
					out<=226;
				end
			end
			1223: begin
				if(in == 0) begin
					state<=1224;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=5122;
					out<=229;
				end
				if(in == 3) begin
					state<=3223;
					out<=230;
				end
				if(in == 4) begin
					state<=7112;
					out<=231;
				end
			end
			1224: begin
				if(in == 0) begin
					state<=1225;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=5123;
					out<=234;
				end
				if(in == 3) begin
					state<=3224;
					out<=235;
				end
				if(in == 4) begin
					state<=7113;
					out<=236;
				end
			end
			1225: begin
				if(in == 0) begin
					state<=1226;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=5124;
					out<=239;
				end
				if(in == 3) begin
					state<=3225;
					out<=240;
				end
				if(in == 4) begin
					state<=7114;
					out<=241;
				end
			end
			1226: begin
				if(in == 0) begin
					state<=1227;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=5125;
					out<=244;
				end
				if(in == 3) begin
					state<=3226;
					out<=245;
				end
				if(in == 4) begin
					state<=7115;
					out<=246;
				end
			end
			1227: begin
				if(in == 0) begin
					state<=1228;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=5126;
					out<=249;
				end
				if(in == 3) begin
					state<=3227;
					out<=250;
				end
				if(in == 4) begin
					state<=7116;
					out<=251;
				end
			end
			1228: begin
				if(in == 0) begin
					state<=1229;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=5127;
					out<=254;
				end
				if(in == 3) begin
					state<=3228;
					out<=255;
				end
				if(in == 4) begin
					state<=7117;
					out<=0;
				end
			end
			1229: begin
				if(in == 0) begin
					state<=1230;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=5128;
					out<=3;
				end
				if(in == 3) begin
					state<=3229;
					out<=4;
				end
				if(in == 4) begin
					state<=7118;
					out<=5;
				end
			end
			1230: begin
				if(in == 0) begin
					state<=691;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=4589;
					out<=8;
				end
				if(in == 3) begin
					state<=2689;
					out<=9;
				end
				if(in == 4) begin
					state<=6578;
					out<=10;
				end
			end
			1231: begin
				if(in == 0) begin
					state<=1232;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=5130;
					out<=13;
				end
				if(in == 3) begin
					state<=2622;
					out<=14;
				end
				if(in == 4) begin
					state<=6511;
					out<=15;
				end
			end
			1232: begin
				if(in == 0) begin
					state<=1233;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=5131;
					out<=18;
				end
				if(in == 3) begin
					state<=2623;
					out<=19;
				end
				if(in == 4) begin
					state<=6512;
					out<=20;
				end
			end
			1233: begin
				if(in == 0) begin
					state<=1234;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=5132;
					out<=23;
				end
				if(in == 3) begin
					state<=2624;
					out<=24;
				end
				if(in == 4) begin
					state<=6513;
					out<=25;
				end
			end
			1234: begin
				if(in == 0) begin
					state<=1235;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=5133;
					out<=28;
				end
				if(in == 3) begin
					state<=2625;
					out<=29;
				end
				if(in == 4) begin
					state<=6514;
					out<=30;
				end
			end
			1235: begin
				if(in == 0) begin
					state<=1236;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=5134;
					out<=33;
				end
				if(in == 3) begin
					state<=2626;
					out<=34;
				end
				if(in == 4) begin
					state<=6515;
					out<=35;
				end
			end
			1236: begin
				if(in == 0) begin
					state<=1237;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=5135;
					out<=38;
				end
				if(in == 3) begin
					state<=2627;
					out<=39;
				end
				if(in == 4) begin
					state<=6516;
					out<=40;
				end
			end
			1237: begin
				if(in == 0) begin
					state<=1238;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=5136;
					out<=43;
				end
				if(in == 3) begin
					state<=2628;
					out<=44;
				end
				if(in == 4) begin
					state<=6517;
					out<=45;
				end
			end
			1238: begin
				if(in == 0) begin
					state<=1239;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=5137;
					out<=48;
				end
				if(in == 3) begin
					state<=2629;
					out<=49;
				end
				if(in == 4) begin
					state<=6518;
					out<=50;
				end
			end
			1239: begin
				if(in == 0) begin
					state<=1240;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=5138;
					out<=53;
				end
				if(in == 3) begin
					state<=2630;
					out<=54;
				end
				if(in == 4) begin
					state<=6519;
					out<=55;
				end
			end
			1240: begin
				if(in == 0) begin
					state<=1241;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=5139;
					out<=58;
				end
				if(in == 3) begin
					state<=2631;
					out<=59;
				end
				if(in == 4) begin
					state<=6520;
					out<=60;
				end
			end
			1241: begin
				if(in == 0) begin
					state<=1242;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=5140;
					out<=63;
				end
				if(in == 3) begin
					state<=2632;
					out<=64;
				end
				if(in == 4) begin
					state<=6521;
					out<=65;
				end
			end
			1242: begin
				if(in == 0) begin
					state<=1243;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=5141;
					out<=68;
				end
				if(in == 3) begin
					state<=2633;
					out<=69;
				end
				if(in == 4) begin
					state<=6522;
					out<=70;
				end
			end
			1243: begin
				if(in == 0) begin
					state<=1244;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=5142;
					out<=73;
				end
				if(in == 3) begin
					state<=2634;
					out<=74;
				end
				if(in == 4) begin
					state<=6523;
					out<=75;
				end
			end
			1244: begin
				if(in == 0) begin
					state<=1245;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=5143;
					out<=78;
				end
				if(in == 3) begin
					state<=2635;
					out<=79;
				end
				if(in == 4) begin
					state<=6524;
					out<=80;
				end
			end
			1245: begin
				if(in == 0) begin
					state<=1246;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=5144;
					out<=83;
				end
				if(in == 3) begin
					state<=2636;
					out<=84;
				end
				if(in == 4) begin
					state<=6525;
					out<=85;
				end
			end
			1246: begin
				if(in == 0) begin
					state<=1247;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=5145;
					out<=88;
				end
				if(in == 3) begin
					state<=2637;
					out<=89;
				end
				if(in == 4) begin
					state<=6526;
					out<=90;
				end
			end
			1247: begin
				if(in == 0) begin
					state<=1248;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=5146;
					out<=93;
				end
				if(in == 3) begin
					state<=2638;
					out<=94;
				end
				if(in == 4) begin
					state<=6527;
					out<=95;
				end
			end
			1248: begin
				if(in == 0) begin
					state<=1249;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=5147;
					out<=98;
				end
				if(in == 3) begin
					state<=2639;
					out<=99;
				end
				if(in == 4) begin
					state<=6528;
					out<=100;
				end
			end
			1249: begin
				if(in == 0) begin
					state<=1250;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=5148;
					out<=103;
				end
				if(in == 3) begin
					state<=2640;
					out<=104;
				end
				if(in == 4) begin
					state<=6529;
					out<=105;
				end
			end
			1250: begin
				if(in == 0) begin
					state<=1251;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=5149;
					out<=108;
				end
				if(in == 3) begin
					state<=2641;
					out<=109;
				end
				if(in == 4) begin
					state<=6530;
					out<=110;
				end
			end
			1251: begin
				if(in == 0) begin
					state<=1252;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=5150;
					out<=113;
				end
				if(in == 3) begin
					state<=2642;
					out<=114;
				end
				if(in == 4) begin
					state<=6531;
					out<=115;
				end
			end
			1252: begin
				if(in == 0) begin
					state<=1253;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=5151;
					out<=118;
				end
				if(in == 3) begin
					state<=2643;
					out<=119;
				end
				if(in == 4) begin
					state<=6532;
					out<=120;
				end
			end
			1253: begin
				if(in == 0) begin
					state<=1254;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=5152;
					out<=123;
				end
				if(in == 3) begin
					state<=2644;
					out<=124;
				end
				if(in == 4) begin
					state<=6533;
					out<=125;
				end
			end
			1254: begin
				if(in == 0) begin
					state<=1255;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=5153;
					out<=128;
				end
				if(in == 3) begin
					state<=2645;
					out<=129;
				end
				if(in == 4) begin
					state<=6534;
					out<=130;
				end
			end
			1255: begin
				if(in == 0) begin
					state<=1256;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=5154;
					out<=133;
				end
				if(in == 3) begin
					state<=2646;
					out<=134;
				end
				if(in == 4) begin
					state<=6535;
					out<=135;
				end
			end
			1256: begin
				if(in == 0) begin
					state<=1257;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=5155;
					out<=138;
				end
				if(in == 3) begin
					state<=2647;
					out<=139;
				end
				if(in == 4) begin
					state<=6536;
					out<=140;
				end
			end
			1257: begin
				if(in == 0) begin
					state<=1258;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=5156;
					out<=143;
				end
				if(in == 3) begin
					state<=2648;
					out<=144;
				end
				if(in == 4) begin
					state<=6537;
					out<=145;
				end
			end
			1258: begin
				if(in == 0) begin
					state<=1259;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=5157;
					out<=148;
				end
				if(in == 3) begin
					state<=2649;
					out<=149;
				end
				if(in == 4) begin
					state<=6538;
					out<=150;
				end
			end
			1259: begin
				if(in == 0) begin
					state<=1260;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=5158;
					out<=153;
				end
				if(in == 3) begin
					state<=2650;
					out<=154;
				end
				if(in == 4) begin
					state<=6539;
					out<=155;
				end
			end
			1260: begin
				if(in == 0) begin
					state<=1261;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=5159;
					out<=158;
				end
				if(in == 3) begin
					state<=2651;
					out<=159;
				end
				if(in == 4) begin
					state<=6540;
					out<=160;
				end
			end
			1261: begin
				if(in == 0) begin
					state<=1262;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=5160;
					out<=163;
				end
				if(in == 3) begin
					state<=2652;
					out<=164;
				end
				if(in == 4) begin
					state<=6541;
					out<=165;
				end
			end
			1262: begin
				if(in == 0) begin
					state<=1263;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=5161;
					out<=168;
				end
				if(in == 3) begin
					state<=2653;
					out<=169;
				end
				if(in == 4) begin
					state<=6542;
					out<=170;
				end
			end
			1263: begin
				if(in == 0) begin
					state<=1264;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=5162;
					out<=173;
				end
				if(in == 3) begin
					state<=2654;
					out<=174;
				end
				if(in == 4) begin
					state<=6543;
					out<=175;
				end
			end
			1264: begin
				if(in == 0) begin
					state<=1265;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=5163;
					out<=178;
				end
				if(in == 3) begin
					state<=2655;
					out<=179;
				end
				if(in == 4) begin
					state<=6544;
					out<=180;
				end
			end
			1265: begin
				if(in == 0) begin
					state<=1266;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=5164;
					out<=183;
				end
				if(in == 3) begin
					state<=2656;
					out<=184;
				end
				if(in == 4) begin
					state<=6545;
					out<=185;
				end
			end
			1266: begin
				if(in == 0) begin
					state<=1267;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=5165;
					out<=188;
				end
				if(in == 3) begin
					state<=2657;
					out<=189;
				end
				if(in == 4) begin
					state<=6546;
					out<=190;
				end
			end
			1267: begin
				if(in == 0) begin
					state<=1268;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=5166;
					out<=193;
				end
				if(in == 3) begin
					state<=2658;
					out<=194;
				end
				if(in == 4) begin
					state<=6547;
					out<=195;
				end
			end
			1268: begin
				if(in == 0) begin
					state<=1269;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=5167;
					out<=198;
				end
				if(in == 3) begin
					state<=2659;
					out<=199;
				end
				if(in == 4) begin
					state<=6548;
					out<=200;
				end
			end
			1269: begin
				if(in == 0) begin
					state<=1270;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=5168;
					out<=203;
				end
				if(in == 3) begin
					state<=2660;
					out<=204;
				end
				if(in == 4) begin
					state<=6549;
					out<=205;
				end
			end
			1270: begin
				if(in == 0) begin
					state<=1271;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=5169;
					out<=208;
				end
				if(in == 3) begin
					state<=2661;
					out<=209;
				end
				if(in == 4) begin
					state<=6550;
					out<=210;
				end
			end
			1271: begin
				if(in == 0) begin
					state<=1272;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=5170;
					out<=213;
				end
				if(in == 3) begin
					state<=2662;
					out<=214;
				end
				if(in == 4) begin
					state<=6551;
					out<=215;
				end
			end
			1272: begin
				if(in == 0) begin
					state<=1273;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=5171;
					out<=218;
				end
				if(in == 3) begin
					state<=2663;
					out<=219;
				end
				if(in == 4) begin
					state<=6552;
					out<=220;
				end
			end
			1273: begin
				if(in == 0) begin
					state<=1274;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=5172;
					out<=223;
				end
				if(in == 3) begin
					state<=2664;
					out<=224;
				end
				if(in == 4) begin
					state<=6553;
					out<=225;
				end
			end
			1274: begin
				if(in == 0) begin
					state<=1275;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=5173;
					out<=228;
				end
				if(in == 3) begin
					state<=2665;
					out<=229;
				end
				if(in == 4) begin
					state<=6554;
					out<=230;
				end
			end
			1275: begin
				if(in == 0) begin
					state<=1276;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=5174;
					out<=233;
				end
				if(in == 3) begin
					state<=2666;
					out<=234;
				end
				if(in == 4) begin
					state<=6555;
					out<=235;
				end
			end
			1276: begin
				if(in == 0) begin
					state<=1277;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=5175;
					out<=238;
				end
				if(in == 3) begin
					state<=2667;
					out<=239;
				end
				if(in == 4) begin
					state<=6556;
					out<=240;
				end
			end
			1277: begin
				if(in == 0) begin
					state<=1278;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=5176;
					out<=243;
				end
				if(in == 3) begin
					state<=2668;
					out<=244;
				end
				if(in == 4) begin
					state<=6557;
					out<=245;
				end
			end
			1278: begin
				if(in == 0) begin
					state<=1279;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=5177;
					out<=248;
				end
				if(in == 3) begin
					state<=2669;
					out<=249;
				end
				if(in == 4) begin
					state<=6558;
					out<=250;
				end
			end
			1279: begin
				if(in == 0) begin
					state<=1280;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=5178;
					out<=253;
				end
				if(in == 3) begin
					state<=3230;
					out<=254;
				end
				if(in == 4) begin
					state<=7119;
					out<=255;
				end
			end
			1280: begin
				if(in == 0) begin
					state<=1281;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=5179;
					out<=2;
				end
				if(in == 3) begin
					state<=3231;
					out<=3;
				end
				if(in == 4) begin
					state<=7120;
					out<=4;
				end
			end
			1281: begin
				if(in == 0) begin
					state<=1282;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=5180;
					out<=7;
				end
				if(in == 3) begin
					state<=3232;
					out<=8;
				end
				if(in == 4) begin
					state<=7121;
					out<=9;
				end
			end
			1282: begin
				if(in == 0) begin
					state<=1283;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=5181;
					out<=12;
				end
				if(in == 3) begin
					state<=3233;
					out<=13;
				end
				if(in == 4) begin
					state<=7122;
					out<=14;
				end
			end
			1283: begin
				if(in == 0) begin
					state<=1284;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=5182;
					out<=17;
				end
				if(in == 3) begin
					state<=3234;
					out<=18;
				end
				if(in == 4) begin
					state<=7123;
					out<=19;
				end
			end
			1284: begin
				if(in == 0) begin
					state<=1285;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=5183;
					out<=22;
				end
				if(in == 3) begin
					state<=3235;
					out<=23;
				end
				if(in == 4) begin
					state<=7124;
					out<=24;
				end
			end
			1285: begin
				if(in == 0) begin
					state<=1286;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=5184;
					out<=27;
				end
				if(in == 3) begin
					state<=3236;
					out<=28;
				end
				if(in == 4) begin
					state<=7125;
					out<=29;
				end
			end
			1286: begin
				if(in == 0) begin
					state<=1287;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=5185;
					out<=32;
				end
				if(in == 3) begin
					state<=3237;
					out<=33;
				end
				if(in == 4) begin
					state<=7126;
					out<=34;
				end
			end
			1287: begin
				if(in == 0) begin
					state<=1288;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=5186;
					out<=37;
				end
				if(in == 3) begin
					state<=3238;
					out<=38;
				end
				if(in == 4) begin
					state<=7127;
					out<=39;
				end
			end
			1288: begin
				if(in == 0) begin
					state<=1289;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=5187;
					out<=42;
				end
				if(in == 3) begin
					state<=3239;
					out<=43;
				end
				if(in == 4) begin
					state<=7128;
					out<=44;
				end
			end
			1289: begin
				if(in == 0) begin
					state<=1290;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=5188;
					out<=47;
				end
				if(in == 3) begin
					state<=3240;
					out<=48;
				end
				if(in == 4) begin
					state<=7129;
					out<=49;
				end
			end
			1290: begin
				if(in == 0) begin
					state<=1291;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=5189;
					out<=52;
				end
				if(in == 3) begin
					state<=3241;
					out<=53;
				end
				if(in == 4) begin
					state<=7130;
					out<=54;
				end
			end
			1291: begin
				if(in == 0) begin
					state<=1292;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=5190;
					out<=57;
				end
				if(in == 3) begin
					state<=3242;
					out<=58;
				end
				if(in == 4) begin
					state<=7131;
					out<=59;
				end
			end
			1292: begin
				if(in == 0) begin
					state<=1293;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=5191;
					out<=62;
				end
				if(in == 3) begin
					state<=3243;
					out<=63;
				end
				if(in == 4) begin
					state<=7132;
					out<=64;
				end
			end
			1293: begin
				if(in == 0) begin
					state<=1294;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=5192;
					out<=67;
				end
				if(in == 3) begin
					state<=3244;
					out<=68;
				end
				if(in == 4) begin
					state<=7133;
					out<=69;
				end
			end
			1294: begin
				if(in == 0) begin
					state<=1295;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=5193;
					out<=72;
				end
				if(in == 3) begin
					state<=3245;
					out<=73;
				end
				if(in == 4) begin
					state<=7134;
					out<=74;
				end
			end
			1295: begin
				if(in == 0) begin
					state<=1296;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=5194;
					out<=77;
				end
				if(in == 3) begin
					state<=3246;
					out<=78;
				end
				if(in == 4) begin
					state<=7135;
					out<=79;
				end
			end
			1296: begin
				if(in == 0) begin
					state<=1297;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=5195;
					out<=82;
				end
				if(in == 3) begin
					state<=3247;
					out<=83;
				end
				if(in == 4) begin
					state<=7136;
					out<=84;
				end
			end
			1297: begin
				if(in == 0) begin
					state<=1298;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=5196;
					out<=87;
				end
				if(in == 3) begin
					state<=3248;
					out<=88;
				end
				if(in == 4) begin
					state<=7137;
					out<=89;
				end
			end
			1298: begin
				if(in == 0) begin
					state<=1299;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=5197;
					out<=92;
				end
				if(in == 3) begin
					state<=3249;
					out<=93;
				end
				if(in == 4) begin
					state<=7138;
					out<=94;
				end
			end
			1299: begin
				if(in == 0) begin
					state<=1300;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=5198;
					out<=97;
				end
				if(in == 3) begin
					state<=3250;
					out<=98;
				end
				if(in == 4) begin
					state<=7139;
					out<=99;
				end
			end
			1300: begin
				if(in == 0) begin
					state<=1301;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=5199;
					out<=102;
				end
				if(in == 3) begin
					state<=3251;
					out<=103;
				end
				if(in == 4) begin
					state<=7140;
					out<=104;
				end
			end
			1301: begin
				if(in == 0) begin
					state<=1302;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=5200;
					out<=107;
				end
				if(in == 3) begin
					state<=3252;
					out<=108;
				end
				if(in == 4) begin
					state<=7141;
					out<=109;
				end
			end
			1302: begin
				if(in == 0) begin
					state<=1303;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=5201;
					out<=112;
				end
				if(in == 3) begin
					state<=3253;
					out<=113;
				end
				if(in == 4) begin
					state<=7142;
					out<=114;
				end
			end
			1303: begin
				if(in == 0) begin
					state<=1304;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=5202;
					out<=117;
				end
				if(in == 3) begin
					state<=3254;
					out<=118;
				end
				if(in == 4) begin
					state<=7143;
					out<=119;
				end
			end
			1304: begin
				if(in == 0) begin
					state<=1305;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=5203;
					out<=122;
				end
				if(in == 3) begin
					state<=3255;
					out<=123;
				end
				if(in == 4) begin
					state<=7144;
					out<=124;
				end
			end
			1305: begin
				if(in == 0) begin
					state<=1306;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=5204;
					out<=127;
				end
				if(in == 3) begin
					state<=3256;
					out<=128;
				end
				if(in == 4) begin
					state<=7145;
					out<=129;
				end
			end
			1306: begin
				if(in == 0) begin
					state<=1307;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=5205;
					out<=132;
				end
				if(in == 3) begin
					state<=3257;
					out<=133;
				end
				if(in == 4) begin
					state<=7146;
					out<=134;
				end
			end
			1307: begin
				if(in == 0) begin
					state<=1308;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=5206;
					out<=137;
				end
				if(in == 3) begin
					state<=3258;
					out<=138;
				end
				if(in == 4) begin
					state<=7147;
					out<=139;
				end
			end
			1308: begin
				if(in == 0) begin
					state<=1309;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=5207;
					out<=142;
				end
				if(in == 3) begin
					state<=3259;
					out<=143;
				end
				if(in == 4) begin
					state<=7148;
					out<=144;
				end
			end
			1309: begin
				if(in == 0) begin
					state<=1310;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=5208;
					out<=147;
				end
				if(in == 3) begin
					state<=3260;
					out<=148;
				end
				if(in == 4) begin
					state<=7149;
					out<=149;
				end
			end
			1310: begin
				if(in == 0) begin
					state<=1311;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=5209;
					out<=152;
				end
				if(in == 3) begin
					state<=2670;
					out<=153;
				end
				if(in == 4) begin
					state<=6559;
					out<=154;
				end
			end
			1311: begin
				if(in == 0) begin
					state<=1312;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=5210;
					out<=157;
				end
				if(in == 3) begin
					state<=2671;
					out<=158;
				end
				if(in == 4) begin
					state<=6560;
					out<=159;
				end
			end
			1312: begin
				if(in == 0) begin
					state<=1313;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=5211;
					out<=162;
				end
				if(in == 3) begin
					state<=2672;
					out<=163;
				end
				if(in == 4) begin
					state<=6561;
					out<=164;
				end
			end
			1313: begin
				if(in == 0) begin
					state<=1314;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=5212;
					out<=167;
				end
				if(in == 3) begin
					state<=2673;
					out<=168;
				end
				if(in == 4) begin
					state<=6562;
					out<=169;
				end
			end
			1314: begin
				if(in == 0) begin
					state<=1315;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=5213;
					out<=172;
				end
				if(in == 3) begin
					state<=2674;
					out<=173;
				end
				if(in == 4) begin
					state<=6563;
					out<=174;
				end
			end
			1315: begin
				if(in == 0) begin
					state<=1316;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=5214;
					out<=177;
				end
				if(in == 3) begin
					state<=2675;
					out<=178;
				end
				if(in == 4) begin
					state<=6564;
					out<=179;
				end
			end
			1316: begin
				if(in == 0) begin
					state<=1317;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=5215;
					out<=182;
				end
				if(in == 3) begin
					state<=2676;
					out<=183;
				end
				if(in == 4) begin
					state<=6565;
					out<=184;
				end
			end
			1317: begin
				if(in == 0) begin
					state<=1318;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=5216;
					out<=187;
				end
				if(in == 3) begin
					state<=2677;
					out<=188;
				end
				if(in == 4) begin
					state<=6566;
					out<=189;
				end
			end
			1318: begin
				if(in == 0) begin
					state<=1319;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=5217;
					out<=192;
				end
				if(in == 3) begin
					state<=2678;
					out<=193;
				end
				if(in == 4) begin
					state<=6567;
					out<=194;
				end
			end
			1319: begin
				if(in == 0) begin
					state<=1320;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=4788;
					out<=197;
				end
				if(in == 3) begin
					state<=2679;
					out<=198;
				end
				if(in == 4) begin
					state<=6568;
					out<=199;
				end
			end
			1320: begin
				if(in == 0) begin
					state<=1321;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=4789;
					out<=202;
				end
				if(in == 3) begin
					state<=2680;
					out<=203;
				end
				if(in == 4) begin
					state<=6569;
					out<=204;
				end
			end
			1321: begin
				if(in == 0) begin
					state<=1322;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=4790;
					out<=207;
				end
				if(in == 3) begin
					state<=2681;
					out<=208;
				end
				if(in == 4) begin
					state<=6570;
					out<=209;
				end
			end
			1322: begin
				if(in == 0) begin
					state<=1323;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=4791;
					out<=212;
				end
				if(in == 3) begin
					state<=2682;
					out<=213;
				end
				if(in == 4) begin
					state<=6571;
					out<=214;
				end
			end
			1323: begin
				if(in == 0) begin
					state<=1324;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=4792;
					out<=217;
				end
				if(in == 3) begin
					state<=2683;
					out<=218;
				end
				if(in == 4) begin
					state<=6572;
					out<=219;
				end
			end
			1324: begin
				if(in == 0) begin
					state<=1325;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=4793;
					out<=222;
				end
				if(in == 3) begin
					state<=2684;
					out<=223;
				end
				if(in == 4) begin
					state<=6573;
					out<=224;
				end
			end
			1325: begin
				if(in == 0) begin
					state<=1326;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=4794;
					out<=227;
				end
				if(in == 3) begin
					state<=2685;
					out<=228;
				end
				if(in == 4) begin
					state<=6574;
					out<=229;
				end
			end
			1326: begin
				if(in == 0) begin
					state<=1327;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=4795;
					out<=232;
				end
				if(in == 3) begin
					state<=2686;
					out<=233;
				end
				if(in == 4) begin
					state<=6575;
					out<=234;
				end
			end
			1327: begin
				if(in == 0) begin
					state<=1328;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=4796;
					out<=237;
				end
				if(in == 3) begin
					state<=2687;
					out<=238;
				end
				if(in == 4) begin
					state<=6576;
					out<=239;
				end
			end
			1328: begin
				if(in == 0) begin
					state<=899;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=4797;
					out<=242;
				end
				if(in == 3) begin
					state<=2688;
					out<=243;
				end
				if(in == 4) begin
					state<=6577;
					out<=244;
				end
			end
			1329: begin
				if(in == 0) begin
					state<=1330;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=5219;
					out<=247;
				end
				if(in == 3) begin
					state<=3262;
					out<=248;
				end
				if(in == 4) begin
					state<=7151;
					out<=249;
				end
			end
			1330: begin
				if(in == 0) begin
					state<=1331;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=5220;
					out<=252;
				end
				if(in == 3) begin
					state<=3263;
					out<=253;
				end
				if(in == 4) begin
					state<=7152;
					out<=254;
				end
			end
			1331: begin
				if(in == 0) begin
					state<=1332;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=5221;
					out<=1;
				end
				if(in == 3) begin
					state<=3264;
					out<=2;
				end
				if(in == 4) begin
					state<=7153;
					out<=3;
				end
			end
			1332: begin
				if(in == 0) begin
					state<=1333;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=5222;
					out<=6;
				end
				if(in == 3) begin
					state<=3265;
					out<=7;
				end
				if(in == 4) begin
					state<=7154;
					out<=8;
				end
			end
			1333: begin
				if(in == 0) begin
					state<=1334;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=5223;
					out<=11;
				end
				if(in == 3) begin
					state<=3266;
					out<=12;
				end
				if(in == 4) begin
					state<=7155;
					out<=13;
				end
			end
			1334: begin
				if(in == 0) begin
					state<=1335;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=5224;
					out<=16;
				end
				if(in == 3) begin
					state<=3267;
					out<=17;
				end
				if(in == 4) begin
					state<=7156;
					out<=18;
				end
			end
			1335: begin
				if(in == 0) begin
					state<=1336;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=5225;
					out<=21;
				end
				if(in == 3) begin
					state<=3268;
					out<=22;
				end
				if(in == 4) begin
					state<=7157;
					out<=23;
				end
			end
			1336: begin
				if(in == 0) begin
					state<=1337;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=5226;
					out<=26;
				end
				if(in == 3) begin
					state<=3269;
					out<=27;
				end
				if(in == 4) begin
					state<=7158;
					out<=28;
				end
			end
			1337: begin
				if(in == 0) begin
					state<=1338;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=5227;
					out<=31;
				end
				if(in == 3) begin
					state<=3270;
					out<=32;
				end
				if(in == 4) begin
					state<=7159;
					out<=33;
				end
			end
			1338: begin
				if(in == 0) begin
					state<=1339;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=5228;
					out<=36;
				end
				if(in == 3) begin
					state<=3271;
					out<=37;
				end
				if(in == 4) begin
					state<=7160;
					out<=38;
				end
			end
			1339: begin
				if(in == 0) begin
					state<=1340;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=5229;
					out<=41;
				end
				if(in == 3) begin
					state<=3272;
					out<=42;
				end
				if(in == 4) begin
					state<=7161;
					out<=43;
				end
			end
			1340: begin
				if(in == 0) begin
					state<=1341;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=5230;
					out<=46;
				end
				if(in == 3) begin
					state<=3273;
					out<=47;
				end
				if(in == 4) begin
					state<=7162;
					out<=48;
				end
			end
			1341: begin
				if(in == 0) begin
					state<=1342;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=5231;
					out<=51;
				end
				if(in == 3) begin
					state<=3274;
					out<=52;
				end
				if(in == 4) begin
					state<=7163;
					out<=53;
				end
			end
			1342: begin
				if(in == 0) begin
					state<=1343;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=5232;
					out<=56;
				end
				if(in == 3) begin
					state<=3275;
					out<=57;
				end
				if(in == 4) begin
					state<=7164;
					out<=58;
				end
			end
			1343: begin
				if(in == 0) begin
					state<=1344;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=5233;
					out<=61;
				end
				if(in == 3) begin
					state<=3276;
					out<=62;
				end
				if(in == 4) begin
					state<=7165;
					out<=63;
				end
			end
			1344: begin
				if(in == 0) begin
					state<=1345;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=5234;
					out<=66;
				end
				if(in == 3) begin
					state<=3277;
					out<=67;
				end
				if(in == 4) begin
					state<=7166;
					out<=68;
				end
			end
			1345: begin
				if(in == 0) begin
					state<=1346;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=5235;
					out<=71;
				end
				if(in == 3) begin
					state<=3278;
					out<=72;
				end
				if(in == 4) begin
					state<=7167;
					out<=73;
				end
			end
			1346: begin
				if(in == 0) begin
					state<=1347;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=5236;
					out<=76;
				end
				if(in == 3) begin
					state<=3279;
					out<=77;
				end
				if(in == 4) begin
					state<=7168;
					out<=78;
				end
			end
			1347: begin
				if(in == 0) begin
					state<=1348;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=5237;
					out<=81;
				end
				if(in == 3) begin
					state<=3280;
					out<=82;
				end
				if(in == 4) begin
					state<=7169;
					out<=83;
				end
			end
			1348: begin
				if(in == 0) begin
					state<=1349;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=5238;
					out<=86;
				end
				if(in == 3) begin
					state<=3281;
					out<=87;
				end
				if(in == 4) begin
					state<=7170;
					out<=88;
				end
			end
			1349: begin
				if(in == 0) begin
					state<=1350;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=5239;
					out<=91;
				end
				if(in == 3) begin
					state<=3282;
					out<=92;
				end
				if(in == 4) begin
					state<=7171;
					out<=93;
				end
			end
			1350: begin
				if(in == 0) begin
					state<=1351;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=5240;
					out<=96;
				end
				if(in == 3) begin
					state<=3283;
					out<=97;
				end
				if(in == 4) begin
					state<=7172;
					out<=98;
				end
			end
			1351: begin
				if(in == 0) begin
					state<=1352;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=5241;
					out<=101;
				end
				if(in == 3) begin
					state<=3284;
					out<=102;
				end
				if(in == 4) begin
					state<=7173;
					out<=103;
				end
			end
			1352: begin
				if(in == 0) begin
					state<=1353;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=5242;
					out<=106;
				end
				if(in == 3) begin
					state<=3285;
					out<=107;
				end
				if(in == 4) begin
					state<=7174;
					out<=108;
				end
			end
			1353: begin
				if(in == 0) begin
					state<=1354;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=5243;
					out<=111;
				end
				if(in == 3) begin
					state<=3286;
					out<=112;
				end
				if(in == 4) begin
					state<=7175;
					out<=113;
				end
			end
			1354: begin
				if(in == 0) begin
					state<=1355;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=5244;
					out<=116;
				end
				if(in == 3) begin
					state<=3287;
					out<=117;
				end
				if(in == 4) begin
					state<=7176;
					out<=118;
				end
			end
			1355: begin
				if(in == 0) begin
					state<=1356;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=5245;
					out<=121;
				end
				if(in == 3) begin
					state<=3288;
					out<=122;
				end
				if(in == 4) begin
					state<=7177;
					out<=123;
				end
			end
			1356: begin
				if(in == 0) begin
					state<=1357;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=5246;
					out<=126;
				end
				if(in == 3) begin
					state<=3289;
					out<=127;
				end
				if(in == 4) begin
					state<=7178;
					out<=128;
				end
			end
			1357: begin
				if(in == 0) begin
					state<=1358;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=5247;
					out<=131;
				end
				if(in == 3) begin
					state<=3290;
					out<=132;
				end
				if(in == 4) begin
					state<=7179;
					out<=133;
				end
			end
			1358: begin
				if(in == 0) begin
					state<=1359;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=5248;
					out<=136;
				end
				if(in == 3) begin
					state<=3291;
					out<=137;
				end
				if(in == 4) begin
					state<=7180;
					out<=138;
				end
			end
			1359: begin
				if(in == 0) begin
					state<=51;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=3949;
					out<=141;
				end
				if(in == 3) begin
					state<=2049;
					out<=142;
				end
				if(in == 4) begin
					state<=5938;
					out<=143;
				end
			end
			1360: begin
				if(in == 0) begin
					state<=1361;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=5250;
					out<=146;
				end
				if(in == 3) begin
					state<=3293;
					out<=147;
				end
				if(in == 4) begin
					state<=7182;
					out<=148;
				end
			end
			1361: begin
				if(in == 0) begin
					state<=1362;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=5251;
					out<=151;
				end
				if(in == 3) begin
					state<=3294;
					out<=152;
				end
				if(in == 4) begin
					state<=7183;
					out<=153;
				end
			end
			1362: begin
				if(in == 0) begin
					state<=1363;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=5252;
					out<=156;
				end
				if(in == 3) begin
					state<=3295;
					out<=157;
				end
				if(in == 4) begin
					state<=7184;
					out<=158;
				end
			end
			1363: begin
				if(in == 0) begin
					state<=1364;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=5253;
					out<=161;
				end
				if(in == 3) begin
					state<=3296;
					out<=162;
				end
				if(in == 4) begin
					state<=7185;
					out<=163;
				end
			end
			1364: begin
				if(in == 0) begin
					state<=1365;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=5254;
					out<=166;
				end
				if(in == 3) begin
					state<=3297;
					out<=167;
				end
				if(in == 4) begin
					state<=7186;
					out<=168;
				end
			end
			1365: begin
				if(in == 0) begin
					state<=1366;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=5255;
					out<=171;
				end
				if(in == 3) begin
					state<=3298;
					out<=172;
				end
				if(in == 4) begin
					state<=7187;
					out<=173;
				end
			end
			1366: begin
				if(in == 0) begin
					state<=1367;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=5256;
					out<=176;
				end
				if(in == 3) begin
					state<=3299;
					out<=177;
				end
				if(in == 4) begin
					state<=7188;
					out<=178;
				end
			end
			1367: begin
				if(in == 0) begin
					state<=1368;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=5257;
					out<=181;
				end
				if(in == 3) begin
					state<=3300;
					out<=182;
				end
				if(in == 4) begin
					state<=7189;
					out<=183;
				end
			end
			1368: begin
				if(in == 0) begin
					state<=1369;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=5258;
					out<=186;
				end
				if(in == 3) begin
					state<=3301;
					out<=187;
				end
				if(in == 4) begin
					state<=7190;
					out<=188;
				end
			end
			1369: begin
				if(in == 0) begin
					state<=1370;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=5259;
					out<=191;
				end
				if(in == 3) begin
					state<=3302;
					out<=192;
				end
				if(in == 4) begin
					state<=7191;
					out<=193;
				end
			end
			1370: begin
				if(in == 0) begin
					state<=1371;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=5260;
					out<=196;
				end
				if(in == 3) begin
					state<=3303;
					out<=197;
				end
				if(in == 4) begin
					state<=7192;
					out<=198;
				end
			end
			1371: begin
				if(in == 0) begin
					state<=1372;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=5261;
					out<=201;
				end
				if(in == 3) begin
					state<=3304;
					out<=202;
				end
				if(in == 4) begin
					state<=7193;
					out<=203;
				end
			end
			1372: begin
				if(in == 0) begin
					state<=1373;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=5262;
					out<=206;
				end
				if(in == 3) begin
					state<=3305;
					out<=207;
				end
				if(in == 4) begin
					state<=7194;
					out<=208;
				end
			end
			1373: begin
				if(in == 0) begin
					state<=1374;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=5263;
					out<=211;
				end
				if(in == 3) begin
					state<=3306;
					out<=212;
				end
				if(in == 4) begin
					state<=7195;
					out<=213;
				end
			end
			1374: begin
				if(in == 0) begin
					state<=1375;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=5264;
					out<=216;
				end
				if(in == 3) begin
					state<=3307;
					out<=217;
				end
				if(in == 4) begin
					state<=7196;
					out<=218;
				end
			end
			1375: begin
				if(in == 0) begin
					state<=1376;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=5265;
					out<=221;
				end
				if(in == 3) begin
					state<=3308;
					out<=222;
				end
				if(in == 4) begin
					state<=7197;
					out<=223;
				end
			end
			1376: begin
				if(in == 0) begin
					state<=1377;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=5266;
					out<=226;
				end
				if(in == 3) begin
					state<=3309;
					out<=227;
				end
				if(in == 4) begin
					state<=7198;
					out<=228;
				end
			end
			1377: begin
				if(in == 0) begin
					state<=1378;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=5267;
					out<=231;
				end
				if(in == 3) begin
					state<=3310;
					out<=232;
				end
				if(in == 4) begin
					state<=7199;
					out<=233;
				end
			end
			1378: begin
				if(in == 0) begin
					state<=1379;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=5268;
					out<=236;
				end
				if(in == 3) begin
					state<=3311;
					out<=237;
				end
				if(in == 4) begin
					state<=7200;
					out<=238;
				end
			end
			1379: begin
				if(in == 0) begin
					state<=1380;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=5269;
					out<=241;
				end
				if(in == 3) begin
					state<=3312;
					out<=242;
				end
				if(in == 4) begin
					state<=7201;
					out<=243;
				end
			end
			1380: begin
				if(in == 0) begin
					state<=1381;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=5270;
					out<=246;
				end
				if(in == 3) begin
					state<=3313;
					out<=247;
				end
				if(in == 4) begin
					state<=7202;
					out<=248;
				end
			end
			1381: begin
				if(in == 0) begin
					state<=1382;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=5271;
					out<=251;
				end
				if(in == 3) begin
					state<=3314;
					out<=252;
				end
				if(in == 4) begin
					state<=7203;
					out<=253;
				end
			end
			1382: begin
				if(in == 0) begin
					state<=1383;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=5272;
					out<=0;
				end
				if(in == 3) begin
					state<=3315;
					out<=1;
				end
				if(in == 4) begin
					state<=7204;
					out<=2;
				end
			end
			1383: begin
				if(in == 0) begin
					state<=1384;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=5273;
					out<=5;
				end
				if(in == 3) begin
					state<=3316;
					out<=6;
				end
				if(in == 4) begin
					state<=7205;
					out<=7;
				end
			end
			1384: begin
				if(in == 0) begin
					state<=1385;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=5274;
					out<=10;
				end
				if(in == 3) begin
					state<=3317;
					out<=11;
				end
				if(in == 4) begin
					state<=7206;
					out<=12;
				end
			end
			1385: begin
				if(in == 0) begin
					state<=1386;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=5275;
					out<=15;
				end
				if(in == 3) begin
					state<=3318;
					out<=16;
				end
				if(in == 4) begin
					state<=7207;
					out<=17;
				end
			end
			1386: begin
				if(in == 0) begin
					state<=1387;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=5276;
					out<=20;
				end
				if(in == 3) begin
					state<=3319;
					out<=21;
				end
				if(in == 4) begin
					state<=7208;
					out<=22;
				end
			end
			1387: begin
				if(in == 0) begin
					state<=1388;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=5277;
					out<=25;
				end
				if(in == 3) begin
					state<=3320;
					out<=26;
				end
				if(in == 4) begin
					state<=7209;
					out<=27;
				end
			end
			1388: begin
				if(in == 0) begin
					state<=1389;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=5278;
					out<=30;
				end
				if(in == 3) begin
					state<=3321;
					out<=31;
				end
				if(in == 4) begin
					state<=7210;
					out<=32;
				end
			end
			1389: begin
				if(in == 0) begin
					state<=1390;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=5279;
					out<=35;
				end
				if(in == 3) begin
					state<=3322;
					out<=36;
				end
				if(in == 4) begin
					state<=7211;
					out<=37;
				end
			end
			1390: begin
				if(in == 0) begin
					state<=120;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=4018;
					out<=40;
				end
				if(in == 3) begin
					state<=2118;
					out<=41;
				end
				if(in == 4) begin
					state<=6007;
					out<=42;
				end
			end
			1391: begin
				if(in == 0) begin
					state<=1392;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=5281;
					out<=45;
				end
				if(in == 3) begin
					state<=3324;
					out<=46;
				end
				if(in == 4) begin
					state<=7213;
					out<=47;
				end
			end
			1392: begin
				if(in == 0) begin
					state<=1393;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=5282;
					out<=50;
				end
				if(in == 3) begin
					state<=3325;
					out<=51;
				end
				if(in == 4) begin
					state<=7214;
					out<=52;
				end
			end
			1393: begin
				if(in == 0) begin
					state<=1394;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=5283;
					out<=55;
				end
				if(in == 3) begin
					state<=3326;
					out<=56;
				end
				if(in == 4) begin
					state<=7215;
					out<=57;
				end
			end
			1394: begin
				if(in == 0) begin
					state<=1395;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=5284;
					out<=60;
				end
				if(in == 3) begin
					state<=3327;
					out<=61;
				end
				if(in == 4) begin
					state<=7216;
					out<=62;
				end
			end
			1395: begin
				if(in == 0) begin
					state<=1396;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=5285;
					out<=65;
				end
				if(in == 3) begin
					state<=3328;
					out<=66;
				end
				if(in == 4) begin
					state<=7217;
					out<=67;
				end
			end
			1396: begin
				if(in == 0) begin
					state<=1397;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=5286;
					out<=70;
				end
				if(in == 3) begin
					state<=3329;
					out<=71;
				end
				if(in == 4) begin
					state<=7218;
					out<=72;
				end
			end
			1397: begin
				if(in == 0) begin
					state<=1398;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=5287;
					out<=75;
				end
				if(in == 3) begin
					state<=3330;
					out<=76;
				end
				if(in == 4) begin
					state<=7219;
					out<=77;
				end
			end
			1398: begin
				if(in == 0) begin
					state<=1399;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=5288;
					out<=80;
				end
				if(in == 3) begin
					state<=3331;
					out<=81;
				end
				if(in == 4) begin
					state<=7220;
					out<=82;
				end
			end
			1399: begin
				if(in == 0) begin
					state<=1400;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=5289;
					out<=85;
				end
				if(in == 3) begin
					state<=3332;
					out<=86;
				end
				if(in == 4) begin
					state<=7221;
					out<=87;
				end
			end
			1400: begin
				if(in == 0) begin
					state<=1401;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=5290;
					out<=90;
				end
				if(in == 3) begin
					state<=3333;
					out<=91;
				end
				if(in == 4) begin
					state<=7222;
					out<=92;
				end
			end
			1401: begin
				if(in == 0) begin
					state<=1402;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=5291;
					out<=95;
				end
				if(in == 3) begin
					state<=3334;
					out<=96;
				end
				if(in == 4) begin
					state<=7223;
					out<=97;
				end
			end
			1402: begin
				if(in == 0) begin
					state<=1403;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=5292;
					out<=100;
				end
				if(in == 3) begin
					state<=3335;
					out<=101;
				end
				if(in == 4) begin
					state<=7224;
					out<=102;
				end
			end
			1403: begin
				if(in == 0) begin
					state<=1404;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=5293;
					out<=105;
				end
				if(in == 3) begin
					state<=3336;
					out<=106;
				end
				if(in == 4) begin
					state<=7225;
					out<=107;
				end
			end
			1404: begin
				if(in == 0) begin
					state<=1405;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=5294;
					out<=110;
				end
				if(in == 3) begin
					state<=3337;
					out<=111;
				end
				if(in == 4) begin
					state<=7226;
					out<=112;
				end
			end
			1405: begin
				if(in == 0) begin
					state<=1406;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=5295;
					out<=115;
				end
				if(in == 3) begin
					state<=3338;
					out<=116;
				end
				if(in == 4) begin
					state<=7227;
					out<=117;
				end
			end
			1406: begin
				if(in == 0) begin
					state<=1407;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=5296;
					out<=120;
				end
				if(in == 3) begin
					state<=3339;
					out<=121;
				end
				if(in == 4) begin
					state<=7228;
					out<=122;
				end
			end
			1407: begin
				if(in == 0) begin
					state<=1408;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=5297;
					out<=125;
				end
				if(in == 3) begin
					state<=3340;
					out<=126;
				end
				if(in == 4) begin
					state<=7229;
					out<=127;
				end
			end
			1408: begin
				if(in == 0) begin
					state<=1409;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=5298;
					out<=130;
				end
				if(in == 3) begin
					state<=3341;
					out<=131;
				end
				if(in == 4) begin
					state<=7230;
					out<=132;
				end
			end
			1409: begin
				if(in == 0) begin
					state<=1410;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=5299;
					out<=135;
				end
				if(in == 3) begin
					state<=3342;
					out<=136;
				end
				if(in == 4) begin
					state<=7231;
					out<=137;
				end
			end
			1410: begin
				if(in == 0) begin
					state<=1411;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=5300;
					out<=140;
				end
				if(in == 3) begin
					state<=3343;
					out<=141;
				end
				if(in == 4) begin
					state<=7232;
					out<=142;
				end
			end
			1411: begin
				if(in == 0) begin
					state<=1412;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=5301;
					out<=145;
				end
				if(in == 3) begin
					state<=3344;
					out<=146;
				end
				if(in == 4) begin
					state<=7233;
					out<=147;
				end
			end
			1412: begin
				if(in == 0) begin
					state<=1413;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=5302;
					out<=150;
				end
				if(in == 3) begin
					state<=3345;
					out<=151;
				end
				if(in == 4) begin
					state<=7234;
					out<=152;
				end
			end
			1413: begin
				if(in == 0) begin
					state<=1414;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=5303;
					out<=155;
				end
				if(in == 3) begin
					state<=3346;
					out<=156;
				end
				if(in == 4) begin
					state<=7235;
					out<=157;
				end
			end
			1414: begin
				if(in == 0) begin
					state<=1415;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=5304;
					out<=160;
				end
				if(in == 3) begin
					state<=3347;
					out<=161;
				end
				if(in == 4) begin
					state<=7236;
					out<=162;
				end
			end
			1415: begin
				if(in == 0) begin
					state<=1416;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=5305;
					out<=165;
				end
				if(in == 3) begin
					state<=3348;
					out<=166;
				end
				if(in == 4) begin
					state<=7237;
					out<=167;
				end
			end
			1416: begin
				if(in == 0) begin
					state<=1417;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=5306;
					out<=170;
				end
				if(in == 3) begin
					state<=3349;
					out<=171;
				end
				if(in == 4) begin
					state<=7238;
					out<=172;
				end
			end
			1417: begin
				if(in == 0) begin
					state<=1418;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=5307;
					out<=175;
				end
				if(in == 3) begin
					state<=3350;
					out<=176;
				end
				if(in == 4) begin
					state<=7239;
					out<=177;
				end
			end
			1418: begin
				if(in == 0) begin
					state<=1419;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=5308;
					out<=180;
				end
				if(in == 3) begin
					state<=3351;
					out<=181;
				end
				if(in == 4) begin
					state<=7240;
					out<=182;
				end
			end
			1419: begin
				if(in == 0) begin
					state<=1420;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=5309;
					out<=185;
				end
				if(in == 3) begin
					state<=3352;
					out<=186;
				end
				if(in == 4) begin
					state<=7241;
					out<=187;
				end
			end
			1420: begin
				if(in == 0) begin
					state<=1421;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=5310;
					out<=190;
				end
				if(in == 3) begin
					state<=3353;
					out<=191;
				end
				if(in == 4) begin
					state<=7242;
					out<=192;
				end
			end
			1421: begin
				if(in == 0) begin
					state<=189;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=4087;
					out<=195;
				end
				if(in == 3) begin
					state<=2187;
					out<=196;
				end
				if(in == 4) begin
					state<=6076;
					out<=197;
				end
			end
			1422: begin
				if(in == 0) begin
					state<=1423;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=5312;
					out<=200;
				end
				if(in == 3) begin
					state<=3355;
					out<=201;
				end
				if(in == 4) begin
					state<=7244;
					out<=202;
				end
			end
			1423: begin
				if(in == 0) begin
					state<=1424;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=5313;
					out<=205;
				end
				if(in == 3) begin
					state<=3356;
					out<=206;
				end
				if(in == 4) begin
					state<=7245;
					out<=207;
				end
			end
			1424: begin
				if(in == 0) begin
					state<=1425;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=5314;
					out<=210;
				end
				if(in == 3) begin
					state<=3357;
					out<=211;
				end
				if(in == 4) begin
					state<=7246;
					out<=212;
				end
			end
			1425: begin
				if(in == 0) begin
					state<=1426;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=5315;
					out<=215;
				end
				if(in == 3) begin
					state<=3358;
					out<=216;
				end
				if(in == 4) begin
					state<=7247;
					out<=217;
				end
			end
			1426: begin
				if(in == 0) begin
					state<=1427;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=5316;
					out<=220;
				end
				if(in == 3) begin
					state<=3359;
					out<=221;
				end
				if(in == 4) begin
					state<=7248;
					out<=222;
				end
			end
			1427: begin
				if(in == 0) begin
					state<=1428;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=5317;
					out<=225;
				end
				if(in == 3) begin
					state<=3360;
					out<=226;
				end
				if(in == 4) begin
					state<=7249;
					out<=227;
				end
			end
			1428: begin
				if(in == 0) begin
					state<=1429;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=5318;
					out<=230;
				end
				if(in == 3) begin
					state<=3361;
					out<=231;
				end
				if(in == 4) begin
					state<=7250;
					out<=232;
				end
			end
			1429: begin
				if(in == 0) begin
					state<=1430;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=5319;
					out<=235;
				end
				if(in == 3) begin
					state<=3362;
					out<=236;
				end
				if(in == 4) begin
					state<=7251;
					out<=237;
				end
			end
			1430: begin
				if(in == 0) begin
					state<=1431;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=5320;
					out<=240;
				end
				if(in == 3) begin
					state<=3363;
					out<=241;
				end
				if(in == 4) begin
					state<=7252;
					out<=242;
				end
			end
			1431: begin
				if(in == 0) begin
					state<=1432;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=5321;
					out<=245;
				end
				if(in == 3) begin
					state<=3364;
					out<=246;
				end
				if(in == 4) begin
					state<=7253;
					out<=247;
				end
			end
			1432: begin
				if(in == 0) begin
					state<=1433;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=5322;
					out<=250;
				end
				if(in == 3) begin
					state<=3365;
					out<=251;
				end
				if(in == 4) begin
					state<=7254;
					out<=252;
				end
			end
			1433: begin
				if(in == 0) begin
					state<=1434;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=5323;
					out<=255;
				end
				if(in == 3) begin
					state<=3366;
					out<=0;
				end
				if(in == 4) begin
					state<=7255;
					out<=1;
				end
			end
			1434: begin
				if(in == 0) begin
					state<=1435;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=5324;
					out<=4;
				end
				if(in == 3) begin
					state<=3367;
					out<=5;
				end
				if(in == 4) begin
					state<=7256;
					out<=6;
				end
			end
			1435: begin
				if(in == 0) begin
					state<=1436;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=5325;
					out<=9;
				end
				if(in == 3) begin
					state<=3368;
					out<=10;
				end
				if(in == 4) begin
					state<=7257;
					out<=11;
				end
			end
			1436: begin
				if(in == 0) begin
					state<=1437;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=5326;
					out<=14;
				end
				if(in == 3) begin
					state<=3369;
					out<=15;
				end
				if(in == 4) begin
					state<=7258;
					out<=16;
				end
			end
			1437: begin
				if(in == 0) begin
					state<=1438;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=5327;
					out<=19;
				end
				if(in == 3) begin
					state<=3370;
					out<=20;
				end
				if(in == 4) begin
					state<=7259;
					out<=21;
				end
			end
			1438: begin
				if(in == 0) begin
					state<=1439;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=5328;
					out<=24;
				end
				if(in == 3) begin
					state<=3371;
					out<=25;
				end
				if(in == 4) begin
					state<=7260;
					out<=26;
				end
			end
			1439: begin
				if(in == 0) begin
					state<=1440;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=5329;
					out<=29;
				end
				if(in == 3) begin
					state<=3372;
					out<=30;
				end
				if(in == 4) begin
					state<=7261;
					out<=31;
				end
			end
			1440: begin
				if(in == 0) begin
					state<=1441;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=5330;
					out<=34;
				end
				if(in == 3) begin
					state<=3373;
					out<=35;
				end
				if(in == 4) begin
					state<=7262;
					out<=36;
				end
			end
			1441: begin
				if(in == 0) begin
					state<=1442;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=5331;
					out<=39;
				end
				if(in == 3) begin
					state<=3374;
					out<=40;
				end
				if(in == 4) begin
					state<=7263;
					out<=41;
				end
			end
			1442: begin
				if(in == 0) begin
					state<=1443;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=5332;
					out<=44;
				end
				if(in == 3) begin
					state<=3375;
					out<=45;
				end
				if(in == 4) begin
					state<=7264;
					out<=46;
				end
			end
			1443: begin
				if(in == 0) begin
					state<=1444;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=5333;
					out<=49;
				end
				if(in == 3) begin
					state<=3376;
					out<=50;
				end
				if(in == 4) begin
					state<=7265;
					out<=51;
				end
			end
			1444: begin
				if(in == 0) begin
					state<=1445;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=5334;
					out<=54;
				end
				if(in == 3) begin
					state<=3377;
					out<=55;
				end
				if(in == 4) begin
					state<=7266;
					out<=56;
				end
			end
			1445: begin
				if(in == 0) begin
					state<=1446;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=5335;
					out<=59;
				end
				if(in == 3) begin
					state<=3378;
					out<=60;
				end
				if(in == 4) begin
					state<=7267;
					out<=61;
				end
			end
			1446: begin
				if(in == 0) begin
					state<=1447;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=5336;
					out<=64;
				end
				if(in == 3) begin
					state<=3379;
					out<=65;
				end
				if(in == 4) begin
					state<=7268;
					out<=66;
				end
			end
			1447: begin
				if(in == 0) begin
					state<=1448;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=5337;
					out<=69;
				end
				if(in == 3) begin
					state<=3380;
					out<=70;
				end
				if(in == 4) begin
					state<=7269;
					out<=71;
				end
			end
			1448: begin
				if(in == 0) begin
					state<=1449;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=5338;
					out<=74;
				end
				if(in == 3) begin
					state<=3381;
					out<=75;
				end
				if(in == 4) begin
					state<=7270;
					out<=76;
				end
			end
			1449: begin
				if(in == 0) begin
					state<=1450;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=5339;
					out<=79;
				end
				if(in == 3) begin
					state<=3382;
					out<=80;
				end
				if(in == 4) begin
					state<=7271;
					out<=81;
				end
			end
			1450: begin
				if(in == 0) begin
					state<=1451;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=5340;
					out<=84;
				end
				if(in == 3) begin
					state<=3383;
					out<=85;
				end
				if(in == 4) begin
					state<=7272;
					out<=86;
				end
			end
			1451: begin
				if(in == 0) begin
					state<=1452;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=5341;
					out<=89;
				end
				if(in == 3) begin
					state<=3384;
					out<=90;
				end
				if(in == 4) begin
					state<=7273;
					out<=91;
				end
			end
			1452: begin
				if(in == 0) begin
					state<=258;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=4156;
					out<=94;
				end
				if(in == 3) begin
					state<=2256;
					out<=95;
				end
				if(in == 4) begin
					state<=6145;
					out<=96;
				end
			end
			1453: begin
				if(in == 0) begin
					state<=1454;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=5343;
					out<=99;
				end
				if(in == 3) begin
					state<=2899;
					out<=100;
				end
				if(in == 4) begin
					state<=6788;
					out<=101;
				end
			end
			1454: begin
				if(in == 0) begin
					state<=1455;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=5344;
					out<=104;
				end
				if(in == 3) begin
					state<=2900;
					out<=105;
				end
				if(in == 4) begin
					state<=6789;
					out<=106;
				end
			end
			1455: begin
				if(in == 0) begin
					state<=1456;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=5345;
					out<=109;
				end
				if(in == 3) begin
					state<=2901;
					out<=110;
				end
				if(in == 4) begin
					state<=6790;
					out<=111;
				end
			end
			1456: begin
				if(in == 0) begin
					state<=1457;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=5346;
					out<=114;
				end
				if(in == 3) begin
					state<=2902;
					out<=115;
				end
				if(in == 4) begin
					state<=6791;
					out<=116;
				end
			end
			1457: begin
				if(in == 0) begin
					state<=1458;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=5347;
					out<=119;
				end
				if(in == 3) begin
					state<=2903;
					out<=120;
				end
				if(in == 4) begin
					state<=6792;
					out<=121;
				end
			end
			1458: begin
				if(in == 0) begin
					state<=1459;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=5348;
					out<=124;
				end
				if(in == 3) begin
					state<=2904;
					out<=125;
				end
				if(in == 4) begin
					state<=6793;
					out<=126;
				end
			end
			1459: begin
				if(in == 0) begin
					state<=1460;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=5349;
					out<=129;
				end
				if(in == 3) begin
					state<=2905;
					out<=130;
				end
				if(in == 4) begin
					state<=6794;
					out<=131;
				end
			end
			1460: begin
				if(in == 0) begin
					state<=1461;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=5350;
					out<=134;
				end
				if(in == 3) begin
					state<=2906;
					out<=135;
				end
				if(in == 4) begin
					state<=6795;
					out<=136;
				end
			end
			1461: begin
				if(in == 0) begin
					state<=1462;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=5351;
					out<=139;
				end
				if(in == 3) begin
					state<=2907;
					out<=140;
				end
				if(in == 4) begin
					state<=6796;
					out<=141;
				end
			end
			1462: begin
				if(in == 0) begin
					state<=1463;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=5352;
					out<=144;
				end
				if(in == 3) begin
					state<=2908;
					out<=145;
				end
				if(in == 4) begin
					state<=6797;
					out<=146;
				end
			end
			1463: begin
				if(in == 0) begin
					state<=1464;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=5353;
					out<=149;
				end
				if(in == 3) begin
					state<=2909;
					out<=150;
				end
				if(in == 4) begin
					state<=6798;
					out<=151;
				end
			end
			1464: begin
				if(in == 0) begin
					state<=1465;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=5354;
					out<=154;
				end
				if(in == 3) begin
					state<=2910;
					out<=155;
				end
				if(in == 4) begin
					state<=6799;
					out<=156;
				end
			end
			1465: begin
				if(in == 0) begin
					state<=1466;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=5355;
					out<=159;
				end
				if(in == 3) begin
					state<=2911;
					out<=160;
				end
				if(in == 4) begin
					state<=6800;
					out<=161;
				end
			end
			1466: begin
				if(in == 0) begin
					state<=1467;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=5356;
					out<=164;
				end
				if(in == 3) begin
					state<=2912;
					out<=165;
				end
				if(in == 4) begin
					state<=6801;
					out<=166;
				end
			end
			1467: begin
				if(in == 0) begin
					state<=1468;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=5357;
					out<=169;
				end
				if(in == 3) begin
					state<=2913;
					out<=170;
				end
				if(in == 4) begin
					state<=6802;
					out<=171;
				end
			end
			1468: begin
				if(in == 0) begin
					state<=1469;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=5358;
					out<=174;
				end
				if(in == 3) begin
					state<=2914;
					out<=175;
				end
				if(in == 4) begin
					state<=6803;
					out<=176;
				end
			end
			1469: begin
				if(in == 0) begin
					state<=1470;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=5359;
					out<=179;
				end
				if(in == 3) begin
					state<=2915;
					out<=180;
				end
				if(in == 4) begin
					state<=6804;
					out<=181;
				end
			end
			1470: begin
				if(in == 0) begin
					state<=1471;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=5360;
					out<=184;
				end
				if(in == 3) begin
					state<=2916;
					out<=185;
				end
				if(in == 4) begin
					state<=6805;
					out<=186;
				end
			end
			1471: begin
				if(in == 0) begin
					state<=1472;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=5361;
					out<=189;
				end
				if(in == 3) begin
					state<=2917;
					out<=190;
				end
				if(in == 4) begin
					state<=6806;
					out<=191;
				end
			end
			1472: begin
				if(in == 0) begin
					state<=1473;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=5362;
					out<=194;
				end
				if(in == 3) begin
					state<=2918;
					out<=195;
				end
				if(in == 4) begin
					state<=6807;
					out<=196;
				end
			end
			1473: begin
				if(in == 0) begin
					state<=1474;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=5363;
					out<=199;
				end
				if(in == 3) begin
					state<=2919;
					out<=200;
				end
				if(in == 4) begin
					state<=6808;
					out<=201;
				end
			end
			1474: begin
				if(in == 0) begin
					state<=1475;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=5364;
					out<=204;
				end
				if(in == 3) begin
					state<=2920;
					out<=205;
				end
				if(in == 4) begin
					state<=6809;
					out<=206;
				end
			end
			1475: begin
				if(in == 0) begin
					state<=1476;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=5365;
					out<=209;
				end
				if(in == 3) begin
					state<=2921;
					out<=210;
				end
				if(in == 4) begin
					state<=6810;
					out<=211;
				end
			end
			1476: begin
				if(in == 0) begin
					state<=1477;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=5366;
					out<=214;
				end
				if(in == 3) begin
					state<=2922;
					out<=215;
				end
				if(in == 4) begin
					state<=6811;
					out<=216;
				end
			end
			1477: begin
				if(in == 0) begin
					state<=1478;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=5367;
					out<=219;
				end
				if(in == 3) begin
					state<=2923;
					out<=220;
				end
				if(in == 4) begin
					state<=6812;
					out<=221;
				end
			end
			1478: begin
				if(in == 0) begin
					state<=1479;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=5368;
					out<=224;
				end
				if(in == 3) begin
					state<=2924;
					out<=225;
				end
				if(in == 4) begin
					state<=6813;
					out<=226;
				end
			end
			1479: begin
				if(in == 0) begin
					state<=1480;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=5369;
					out<=229;
				end
				if(in == 3) begin
					state<=2925;
					out<=230;
				end
				if(in == 4) begin
					state<=6814;
					out<=231;
				end
			end
			1480: begin
				if(in == 0) begin
					state<=1481;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=5370;
					out<=234;
				end
				if(in == 3) begin
					state<=2926;
					out<=235;
				end
				if(in == 4) begin
					state<=6815;
					out<=236;
				end
			end
			1481: begin
				if(in == 0) begin
					state<=1482;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=5371;
					out<=239;
				end
				if(in == 3) begin
					state<=2927;
					out<=240;
				end
				if(in == 4) begin
					state<=6816;
					out<=241;
				end
			end
			1482: begin
				if(in == 0) begin
					state<=1483;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=5372;
					out<=244;
				end
				if(in == 3) begin
					state<=2928;
					out<=245;
				end
				if(in == 4) begin
					state<=6817;
					out<=246;
				end
			end
			1483: begin
				if(in == 0) begin
					state<=327;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=4225;
					out<=249;
				end
				if(in == 3) begin
					state<=2325;
					out<=250;
				end
				if(in == 4) begin
					state<=6214;
					out<=251;
				end
			end
			1484: begin
				if(in == 0) begin
					state<=1485;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=5374;
					out<=254;
				end
				if(in == 3) begin
					state<=3417;
					out<=255;
				end
				if(in == 4) begin
					state<=7306;
					out<=0;
				end
			end
			1485: begin
				if(in == 0) begin
					state<=1486;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=5375;
					out<=3;
				end
				if(in == 3) begin
					state<=3418;
					out<=4;
				end
				if(in == 4) begin
					state<=7307;
					out<=5;
				end
			end
			1486: begin
				if(in == 0) begin
					state<=1487;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=5376;
					out<=8;
				end
				if(in == 3) begin
					state<=3419;
					out<=9;
				end
				if(in == 4) begin
					state<=7308;
					out<=10;
				end
			end
			1487: begin
				if(in == 0) begin
					state<=1488;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=5377;
					out<=13;
				end
				if(in == 3) begin
					state<=3420;
					out<=14;
				end
				if(in == 4) begin
					state<=7309;
					out<=15;
				end
			end
			1488: begin
				if(in == 0) begin
					state<=1489;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=5378;
					out<=18;
				end
				if(in == 3) begin
					state<=3421;
					out<=19;
				end
				if(in == 4) begin
					state<=7310;
					out<=20;
				end
			end
			1489: begin
				if(in == 0) begin
					state<=1490;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=5379;
					out<=23;
				end
				if(in == 3) begin
					state<=3422;
					out<=24;
				end
				if(in == 4) begin
					state<=7311;
					out<=25;
				end
			end
			1490: begin
				if(in == 0) begin
					state<=1491;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=5380;
					out<=28;
				end
				if(in == 3) begin
					state<=3423;
					out<=29;
				end
				if(in == 4) begin
					state<=7312;
					out<=30;
				end
			end
			1491: begin
				if(in == 0) begin
					state<=1492;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=5381;
					out<=33;
				end
				if(in == 3) begin
					state<=3424;
					out<=34;
				end
				if(in == 4) begin
					state<=7313;
					out<=35;
				end
			end
			1492: begin
				if(in == 0) begin
					state<=1493;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=5382;
					out<=38;
				end
				if(in == 3) begin
					state<=3425;
					out<=39;
				end
				if(in == 4) begin
					state<=7314;
					out<=40;
				end
			end
			1493: begin
				if(in == 0) begin
					state<=1494;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=5383;
					out<=43;
				end
				if(in == 3) begin
					state<=3426;
					out<=44;
				end
				if(in == 4) begin
					state<=7315;
					out<=45;
				end
			end
			1494: begin
				if(in == 0) begin
					state<=1495;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=5384;
					out<=48;
				end
				if(in == 3) begin
					state<=3427;
					out<=49;
				end
				if(in == 4) begin
					state<=7316;
					out<=50;
				end
			end
			1495: begin
				if(in == 0) begin
					state<=1496;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=5385;
					out<=53;
				end
				if(in == 3) begin
					state<=3428;
					out<=54;
				end
				if(in == 4) begin
					state<=7317;
					out<=55;
				end
			end
			1496: begin
				if(in == 0) begin
					state<=1497;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=5386;
					out<=58;
				end
				if(in == 3) begin
					state<=3429;
					out<=59;
				end
				if(in == 4) begin
					state<=7318;
					out<=60;
				end
			end
			1497: begin
				if(in == 0) begin
					state<=1498;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=5387;
					out<=63;
				end
				if(in == 3) begin
					state<=3430;
					out<=64;
				end
				if(in == 4) begin
					state<=7319;
					out<=65;
				end
			end
			1498: begin
				if(in == 0) begin
					state<=1499;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=5388;
					out<=68;
				end
				if(in == 3) begin
					state<=3431;
					out<=69;
				end
				if(in == 4) begin
					state<=7320;
					out<=70;
				end
			end
			1499: begin
				if(in == 0) begin
					state<=1500;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=5389;
					out<=73;
				end
				if(in == 3) begin
					state<=3432;
					out<=74;
				end
				if(in == 4) begin
					state<=7321;
					out<=75;
				end
			end
			1500: begin
				if(in == 0) begin
					state<=1501;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=5390;
					out<=78;
				end
				if(in == 3) begin
					state<=3433;
					out<=79;
				end
				if(in == 4) begin
					state<=7322;
					out<=80;
				end
			end
			1501: begin
				if(in == 0) begin
					state<=1502;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=5391;
					out<=83;
				end
				if(in == 3) begin
					state<=3434;
					out<=84;
				end
				if(in == 4) begin
					state<=7323;
					out<=85;
				end
			end
			1502: begin
				if(in == 0) begin
					state<=1503;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=5392;
					out<=88;
				end
				if(in == 3) begin
					state<=3435;
					out<=89;
				end
				if(in == 4) begin
					state<=7324;
					out<=90;
				end
			end
			1503: begin
				if(in == 0) begin
					state<=1504;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=5393;
					out<=93;
				end
				if(in == 3) begin
					state<=3436;
					out<=94;
				end
				if(in == 4) begin
					state<=7325;
					out<=95;
				end
			end
			1504: begin
				if(in == 0) begin
					state<=1505;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=5394;
					out<=98;
				end
				if(in == 3) begin
					state<=3437;
					out<=99;
				end
				if(in == 4) begin
					state<=7326;
					out<=100;
				end
			end
			1505: begin
				if(in == 0) begin
					state<=1506;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=5395;
					out<=103;
				end
				if(in == 3) begin
					state<=3438;
					out<=104;
				end
				if(in == 4) begin
					state<=7327;
					out<=105;
				end
			end
			1506: begin
				if(in == 0) begin
					state<=1507;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=5396;
					out<=108;
				end
				if(in == 3) begin
					state<=3439;
					out<=109;
				end
				if(in == 4) begin
					state<=7328;
					out<=110;
				end
			end
			1507: begin
				if(in == 0) begin
					state<=1508;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=5397;
					out<=113;
				end
				if(in == 3) begin
					state<=3440;
					out<=114;
				end
				if(in == 4) begin
					state<=7329;
					out<=115;
				end
			end
			1508: begin
				if(in == 0) begin
					state<=1509;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=5398;
					out<=118;
				end
				if(in == 3) begin
					state<=3441;
					out<=119;
				end
				if(in == 4) begin
					state<=7330;
					out<=120;
				end
			end
			1509: begin
				if(in == 0) begin
					state<=1510;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=5399;
					out<=123;
				end
				if(in == 3) begin
					state<=3442;
					out<=124;
				end
				if(in == 4) begin
					state<=7331;
					out<=125;
				end
			end
			1510: begin
				if(in == 0) begin
					state<=1511;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=5400;
					out<=128;
				end
				if(in == 3) begin
					state<=3443;
					out<=129;
				end
				if(in == 4) begin
					state<=7332;
					out<=130;
				end
			end
			1511: begin
				if(in == 0) begin
					state<=1512;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=5401;
					out<=133;
				end
				if(in == 3) begin
					state<=3444;
					out<=134;
				end
				if(in == 4) begin
					state<=7333;
					out<=135;
				end
			end
			1512: begin
				if(in == 0) begin
					state<=1513;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=5402;
					out<=138;
				end
				if(in == 3) begin
					state<=3445;
					out<=139;
				end
				if(in == 4) begin
					state<=7334;
					out<=140;
				end
			end
			1513: begin
				if(in == 0) begin
					state<=1514;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=5403;
					out<=143;
				end
				if(in == 3) begin
					state<=3446;
					out<=144;
				end
				if(in == 4) begin
					state<=7335;
					out<=145;
				end
			end
			1514: begin
				if(in == 0) begin
					state<=465;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=4363;
					out<=148;
				end
				if(in == 3) begin
					state<=2463;
					out<=149;
				end
				if(in == 4) begin
					state<=6352;
					out<=150;
				end
			end
			1515: begin
				if(in == 0) begin
					state<=1516;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=5405;
					out<=153;
				end
				if(in == 3) begin
					state<=3448;
					out<=154;
				end
				if(in == 4) begin
					state<=7337;
					out<=155;
				end
			end
			1516: begin
				if(in == 0) begin
					state<=1517;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=5406;
					out<=158;
				end
				if(in == 3) begin
					state<=3449;
					out<=159;
				end
				if(in == 4) begin
					state<=7338;
					out<=160;
				end
			end
			1517: begin
				if(in == 0) begin
					state<=1518;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=5407;
					out<=163;
				end
				if(in == 3) begin
					state<=3450;
					out<=164;
				end
				if(in == 4) begin
					state<=7339;
					out<=165;
				end
			end
			1518: begin
				if(in == 0) begin
					state<=1519;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=5408;
					out<=168;
				end
				if(in == 3) begin
					state<=3451;
					out<=169;
				end
				if(in == 4) begin
					state<=7340;
					out<=170;
				end
			end
			1519: begin
				if(in == 0) begin
					state<=1520;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=5409;
					out<=173;
				end
				if(in == 3) begin
					state<=3452;
					out<=174;
				end
				if(in == 4) begin
					state<=7341;
					out<=175;
				end
			end
			1520: begin
				if(in == 0) begin
					state<=1521;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=5410;
					out<=178;
				end
				if(in == 3) begin
					state<=3453;
					out<=179;
				end
				if(in == 4) begin
					state<=7342;
					out<=180;
				end
			end
			1521: begin
				if(in == 0) begin
					state<=1522;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=5411;
					out<=183;
				end
				if(in == 3) begin
					state<=3454;
					out<=184;
				end
				if(in == 4) begin
					state<=7343;
					out<=185;
				end
			end
			1522: begin
				if(in == 0) begin
					state<=1523;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=5412;
					out<=188;
				end
				if(in == 3) begin
					state<=3455;
					out<=189;
				end
				if(in == 4) begin
					state<=7344;
					out<=190;
				end
			end
			1523: begin
				if(in == 0) begin
					state<=1524;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=5413;
					out<=193;
				end
				if(in == 3) begin
					state<=3456;
					out<=194;
				end
				if(in == 4) begin
					state<=7345;
					out<=195;
				end
			end
			1524: begin
				if(in == 0) begin
					state<=1525;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=5414;
					out<=198;
				end
				if(in == 3) begin
					state<=3457;
					out<=199;
				end
				if(in == 4) begin
					state<=7346;
					out<=200;
				end
			end
			1525: begin
				if(in == 0) begin
					state<=1526;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=5415;
					out<=203;
				end
				if(in == 3) begin
					state<=3458;
					out<=204;
				end
				if(in == 4) begin
					state<=7347;
					out<=205;
				end
			end
			1526: begin
				if(in == 0) begin
					state<=1527;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=5416;
					out<=208;
				end
				if(in == 3) begin
					state<=3459;
					out<=209;
				end
				if(in == 4) begin
					state<=7348;
					out<=210;
				end
			end
			1527: begin
				if(in == 0) begin
					state<=1528;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=5417;
					out<=213;
				end
				if(in == 3) begin
					state<=3460;
					out<=214;
				end
				if(in == 4) begin
					state<=7349;
					out<=215;
				end
			end
			1528: begin
				if(in == 0) begin
					state<=1529;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=5418;
					out<=218;
				end
				if(in == 3) begin
					state<=3461;
					out<=219;
				end
				if(in == 4) begin
					state<=7350;
					out<=220;
				end
			end
			1529: begin
				if(in == 0) begin
					state<=1530;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=5419;
					out<=223;
				end
				if(in == 3) begin
					state<=3462;
					out<=224;
				end
				if(in == 4) begin
					state<=7351;
					out<=225;
				end
			end
			1530: begin
				if(in == 0) begin
					state<=1531;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=5420;
					out<=228;
				end
				if(in == 3) begin
					state<=3463;
					out<=229;
				end
				if(in == 4) begin
					state<=7352;
					out<=230;
				end
			end
			1531: begin
				if(in == 0) begin
					state<=1532;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=5421;
					out<=233;
				end
				if(in == 3) begin
					state<=3464;
					out<=234;
				end
				if(in == 4) begin
					state<=7353;
					out<=235;
				end
			end
			1532: begin
				if(in == 0) begin
					state<=1533;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=5422;
					out<=238;
				end
				if(in == 3) begin
					state<=3465;
					out<=239;
				end
				if(in == 4) begin
					state<=7354;
					out<=240;
				end
			end
			1533: begin
				if(in == 0) begin
					state<=1534;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=5423;
					out<=243;
				end
				if(in == 3) begin
					state<=3466;
					out<=244;
				end
				if(in == 4) begin
					state<=7355;
					out<=245;
				end
			end
			1534: begin
				if(in == 0) begin
					state<=1535;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=5424;
					out<=248;
				end
				if(in == 3) begin
					state<=3467;
					out<=249;
				end
				if(in == 4) begin
					state<=7356;
					out<=250;
				end
			end
			1535: begin
				if(in == 0) begin
					state<=1536;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=5425;
					out<=253;
				end
				if(in == 3) begin
					state<=3468;
					out<=254;
				end
				if(in == 4) begin
					state<=7357;
					out<=255;
				end
			end
			1536: begin
				if(in == 0) begin
					state<=1537;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=5426;
					out<=2;
				end
				if(in == 3) begin
					state<=3469;
					out<=3;
				end
				if(in == 4) begin
					state<=7358;
					out<=4;
				end
			end
			1537: begin
				if(in == 0) begin
					state<=1538;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=5427;
					out<=7;
				end
				if(in == 3) begin
					state<=3470;
					out<=8;
				end
				if(in == 4) begin
					state<=7359;
					out<=9;
				end
			end
			1538: begin
				if(in == 0) begin
					state<=1539;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=5428;
					out<=12;
				end
				if(in == 3) begin
					state<=3471;
					out<=13;
				end
				if(in == 4) begin
					state<=7360;
					out<=14;
				end
			end
			1539: begin
				if(in == 0) begin
					state<=1540;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=5429;
					out<=17;
				end
				if(in == 3) begin
					state<=3472;
					out<=18;
				end
				if(in == 4) begin
					state<=7361;
					out<=19;
				end
			end
			1540: begin
				if(in == 0) begin
					state<=1541;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=5430;
					out<=22;
				end
				if(in == 3) begin
					state<=3473;
					out<=23;
				end
				if(in == 4) begin
					state<=7362;
					out<=24;
				end
			end
			1541: begin
				if(in == 0) begin
					state<=1542;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=5431;
					out<=27;
				end
				if(in == 3) begin
					state<=3474;
					out<=28;
				end
				if(in == 4) begin
					state<=7363;
					out<=29;
				end
			end
			1542: begin
				if(in == 0) begin
					state<=1543;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=5432;
					out<=32;
				end
				if(in == 3) begin
					state<=3475;
					out<=33;
				end
				if(in == 4) begin
					state<=7364;
					out<=34;
				end
			end
			1543: begin
				if(in == 0) begin
					state<=1544;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=5433;
					out<=37;
				end
				if(in == 3) begin
					state<=3476;
					out<=38;
				end
				if(in == 4) begin
					state<=7365;
					out<=39;
				end
			end
			1544: begin
				if(in == 0) begin
					state<=1545;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=5434;
					out<=42;
				end
				if(in == 3) begin
					state<=3477;
					out<=43;
				end
				if(in == 4) begin
					state<=7366;
					out<=44;
				end
			end
			1545: begin
				if(in == 0) begin
					state<=534;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=4432;
					out<=47;
				end
				if(in == 3) begin
					state<=2532;
					out<=48;
				end
				if(in == 4) begin
					state<=6421;
					out<=49;
				end
			end
			1546: begin
				if(in == 0) begin
					state<=1547;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=5436;
					out<=52;
				end
				if(in == 3) begin
					state<=3479;
					out<=53;
				end
				if(in == 4) begin
					state<=7368;
					out<=54;
				end
			end
			1547: begin
				if(in == 0) begin
					state<=1548;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=5437;
					out<=57;
				end
				if(in == 3) begin
					state<=3480;
					out<=58;
				end
				if(in == 4) begin
					state<=7369;
					out<=59;
				end
			end
			1548: begin
				if(in == 0) begin
					state<=1549;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=5438;
					out<=62;
				end
				if(in == 3) begin
					state<=3481;
					out<=63;
				end
				if(in == 4) begin
					state<=7370;
					out<=64;
				end
			end
			1549: begin
				if(in == 0) begin
					state<=1550;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=5439;
					out<=67;
				end
				if(in == 3) begin
					state<=3482;
					out<=68;
				end
				if(in == 4) begin
					state<=7371;
					out<=69;
				end
			end
			1550: begin
				if(in == 0) begin
					state<=1551;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=5440;
					out<=72;
				end
				if(in == 3) begin
					state<=3483;
					out<=73;
				end
				if(in == 4) begin
					state<=7372;
					out<=74;
				end
			end
			1551: begin
				if(in == 0) begin
					state<=1552;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=5441;
					out<=77;
				end
				if(in == 3) begin
					state<=3484;
					out<=78;
				end
				if(in == 4) begin
					state<=7373;
					out<=79;
				end
			end
			1552: begin
				if(in == 0) begin
					state<=1553;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=5442;
					out<=82;
				end
				if(in == 3) begin
					state<=3485;
					out<=83;
				end
				if(in == 4) begin
					state<=7374;
					out<=84;
				end
			end
			1553: begin
				if(in == 0) begin
					state<=1554;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=5443;
					out<=87;
				end
				if(in == 3) begin
					state<=3486;
					out<=88;
				end
				if(in == 4) begin
					state<=7375;
					out<=89;
				end
			end
			1554: begin
				if(in == 0) begin
					state<=1555;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=5444;
					out<=92;
				end
				if(in == 3) begin
					state<=3487;
					out<=93;
				end
				if(in == 4) begin
					state<=7376;
					out<=94;
				end
			end
			1555: begin
				if(in == 0) begin
					state<=1556;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=5445;
					out<=97;
				end
				if(in == 3) begin
					state<=3488;
					out<=98;
				end
				if(in == 4) begin
					state<=7377;
					out<=99;
				end
			end
			1556: begin
				if(in == 0) begin
					state<=1557;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=5446;
					out<=102;
				end
				if(in == 3) begin
					state<=3489;
					out<=103;
				end
				if(in == 4) begin
					state<=7378;
					out<=104;
				end
			end
			1557: begin
				if(in == 0) begin
					state<=1558;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=5447;
					out<=107;
				end
				if(in == 3) begin
					state<=3490;
					out<=108;
				end
				if(in == 4) begin
					state<=7379;
					out<=109;
				end
			end
			1558: begin
				if(in == 0) begin
					state<=1559;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=5448;
					out<=112;
				end
				if(in == 3) begin
					state<=3491;
					out<=113;
				end
				if(in == 4) begin
					state<=7380;
					out<=114;
				end
			end
			1559: begin
				if(in == 0) begin
					state<=1560;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=5449;
					out<=117;
				end
				if(in == 3) begin
					state<=3492;
					out<=118;
				end
				if(in == 4) begin
					state<=7381;
					out<=119;
				end
			end
			1560: begin
				if(in == 0) begin
					state<=1561;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=5450;
					out<=122;
				end
				if(in == 3) begin
					state<=3493;
					out<=123;
				end
				if(in == 4) begin
					state<=7382;
					out<=124;
				end
			end
			1561: begin
				if(in == 0) begin
					state<=1562;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=5451;
					out<=127;
				end
				if(in == 3) begin
					state<=3494;
					out<=128;
				end
				if(in == 4) begin
					state<=7383;
					out<=129;
				end
			end
			1562: begin
				if(in == 0) begin
					state<=1563;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=5452;
					out<=132;
				end
				if(in == 3) begin
					state<=3495;
					out<=133;
				end
				if(in == 4) begin
					state<=7384;
					out<=134;
				end
			end
			1563: begin
				if(in == 0) begin
					state<=1564;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=5453;
					out<=137;
				end
				if(in == 3) begin
					state<=3496;
					out<=138;
				end
				if(in == 4) begin
					state<=7385;
					out<=139;
				end
			end
			1564: begin
				if(in == 0) begin
					state<=1565;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=5454;
					out<=142;
				end
				if(in == 3) begin
					state<=3497;
					out<=143;
				end
				if(in == 4) begin
					state<=7386;
					out<=144;
				end
			end
			1565: begin
				if(in == 0) begin
					state<=1566;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=5455;
					out<=147;
				end
				if(in == 3) begin
					state<=3498;
					out<=148;
				end
				if(in == 4) begin
					state<=7387;
					out<=149;
				end
			end
			1566: begin
				if(in == 0) begin
					state<=1567;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=5456;
					out<=152;
				end
				if(in == 3) begin
					state<=3499;
					out<=153;
				end
				if(in == 4) begin
					state<=7388;
					out<=154;
				end
			end
			1567: begin
				if(in == 0) begin
					state<=1568;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=5457;
					out<=157;
				end
				if(in == 3) begin
					state<=3500;
					out<=158;
				end
				if(in == 4) begin
					state<=7389;
					out<=159;
				end
			end
			1568: begin
				if(in == 0) begin
					state<=1569;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=5458;
					out<=162;
				end
				if(in == 3) begin
					state<=3501;
					out<=163;
				end
				if(in == 4) begin
					state<=7390;
					out<=164;
				end
			end
			1569: begin
				if(in == 0) begin
					state<=1570;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=5459;
					out<=167;
				end
				if(in == 3) begin
					state<=3502;
					out<=168;
				end
				if(in == 4) begin
					state<=7391;
					out<=169;
				end
			end
			1570: begin
				if(in == 0) begin
					state<=1571;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=5460;
					out<=172;
				end
				if(in == 3) begin
					state<=3503;
					out<=173;
				end
				if(in == 4) begin
					state<=7392;
					out<=174;
				end
			end
			1571: begin
				if(in == 0) begin
					state<=1572;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=5461;
					out<=177;
				end
				if(in == 3) begin
					state<=3504;
					out<=178;
				end
				if(in == 4) begin
					state<=7393;
					out<=179;
				end
			end
			1572: begin
				if(in == 0) begin
					state<=1573;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=5462;
					out<=182;
				end
				if(in == 3) begin
					state<=3505;
					out<=183;
				end
				if(in == 4) begin
					state<=7394;
					out<=184;
				end
			end
			1573: begin
				if(in == 0) begin
					state<=1574;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=5463;
					out<=187;
				end
				if(in == 3) begin
					state<=3506;
					out<=188;
				end
				if(in == 4) begin
					state<=7395;
					out<=189;
				end
			end
			1574: begin
				if(in == 0) begin
					state<=1575;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=5464;
					out<=192;
				end
				if(in == 3) begin
					state<=3507;
					out<=193;
				end
				if(in == 4) begin
					state<=7396;
					out<=194;
				end
			end
			1575: begin
				if(in == 0) begin
					state<=1576;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=5465;
					out<=197;
				end
				if(in == 3) begin
					state<=3508;
					out<=198;
				end
				if(in == 4) begin
					state<=7397;
					out<=199;
				end
			end
			1576: begin
				if(in == 0) begin
					state<=603;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=4501;
					out<=202;
				end
				if(in == 3) begin
					state<=2601;
					out<=203;
				end
				if(in == 4) begin
					state<=6490;
					out<=204;
				end
			end
			1577: begin
				if(in == 0) begin
					state<=1578;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=5467;
					out<=207;
				end
				if(in == 3) begin
					state<=3231;
					out<=208;
				end
				if(in == 4) begin
					state<=7120;
					out<=209;
				end
			end
			1578: begin
				if(in == 0) begin
					state<=1579;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=5468;
					out<=212;
				end
				if(in == 3) begin
					state<=3232;
					out<=213;
				end
				if(in == 4) begin
					state<=7121;
					out<=214;
				end
			end
			1579: begin
				if(in == 0) begin
					state<=1580;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=5469;
					out<=217;
				end
				if(in == 3) begin
					state<=3233;
					out<=218;
				end
				if(in == 4) begin
					state<=7122;
					out<=219;
				end
			end
			1580: begin
				if(in == 0) begin
					state<=1581;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=5470;
					out<=222;
				end
				if(in == 3) begin
					state<=3234;
					out<=223;
				end
				if(in == 4) begin
					state<=7123;
					out<=224;
				end
			end
			1581: begin
				if(in == 0) begin
					state<=1582;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=5471;
					out<=227;
				end
				if(in == 3) begin
					state<=3235;
					out<=228;
				end
				if(in == 4) begin
					state<=7124;
					out<=229;
				end
			end
			1582: begin
				if(in == 0) begin
					state<=1583;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=5472;
					out<=232;
				end
				if(in == 3) begin
					state<=3236;
					out<=233;
				end
				if(in == 4) begin
					state<=7125;
					out<=234;
				end
			end
			1583: begin
				if(in == 0) begin
					state<=1584;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=5473;
					out<=237;
				end
				if(in == 3) begin
					state<=3237;
					out<=238;
				end
				if(in == 4) begin
					state<=7126;
					out<=239;
				end
			end
			1584: begin
				if(in == 0) begin
					state<=1585;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=5474;
					out<=242;
				end
				if(in == 3) begin
					state<=3238;
					out<=243;
				end
				if(in == 4) begin
					state<=7127;
					out<=244;
				end
			end
			1585: begin
				if(in == 0) begin
					state<=1586;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=5475;
					out<=247;
				end
				if(in == 3) begin
					state<=3239;
					out<=248;
				end
				if(in == 4) begin
					state<=7128;
					out<=249;
				end
			end
			1586: begin
				if(in == 0) begin
					state<=1587;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=5476;
					out<=252;
				end
				if(in == 3) begin
					state<=3240;
					out<=253;
				end
				if(in == 4) begin
					state<=7129;
					out<=254;
				end
			end
			1587: begin
				if(in == 0) begin
					state<=1588;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=5477;
					out<=1;
				end
				if(in == 3) begin
					state<=3241;
					out<=2;
				end
				if(in == 4) begin
					state<=7130;
					out<=3;
				end
			end
			1588: begin
				if(in == 0) begin
					state<=1589;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=5478;
					out<=6;
				end
				if(in == 3) begin
					state<=3242;
					out<=7;
				end
				if(in == 4) begin
					state<=7131;
					out<=8;
				end
			end
			1589: begin
				if(in == 0) begin
					state<=1590;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=5479;
					out<=11;
				end
				if(in == 3) begin
					state<=3243;
					out<=12;
				end
				if(in == 4) begin
					state<=7132;
					out<=13;
				end
			end
			1590: begin
				if(in == 0) begin
					state<=1591;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=5480;
					out<=16;
				end
				if(in == 3) begin
					state<=3244;
					out<=17;
				end
				if(in == 4) begin
					state<=7133;
					out<=18;
				end
			end
			1591: begin
				if(in == 0) begin
					state<=1592;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=5481;
					out<=21;
				end
				if(in == 3) begin
					state<=3245;
					out<=22;
				end
				if(in == 4) begin
					state<=7134;
					out<=23;
				end
			end
			1592: begin
				if(in == 0) begin
					state<=1593;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=5482;
					out<=26;
				end
				if(in == 3) begin
					state<=3246;
					out<=27;
				end
				if(in == 4) begin
					state<=7135;
					out<=28;
				end
			end
			1593: begin
				if(in == 0) begin
					state<=1594;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=5483;
					out<=31;
				end
				if(in == 3) begin
					state<=3247;
					out<=32;
				end
				if(in == 4) begin
					state<=7136;
					out<=33;
				end
			end
			1594: begin
				if(in == 0) begin
					state<=1595;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=5484;
					out<=36;
				end
				if(in == 3) begin
					state<=3248;
					out<=37;
				end
				if(in == 4) begin
					state<=7137;
					out<=38;
				end
			end
			1595: begin
				if(in == 0) begin
					state<=1596;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=5485;
					out<=41;
				end
				if(in == 3) begin
					state<=3249;
					out<=42;
				end
				if(in == 4) begin
					state<=7138;
					out<=43;
				end
			end
			1596: begin
				if(in == 0) begin
					state<=1597;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=5486;
					out<=46;
				end
				if(in == 3) begin
					state<=3250;
					out<=47;
				end
				if(in == 4) begin
					state<=7139;
					out<=48;
				end
			end
			1597: begin
				if(in == 0) begin
					state<=1598;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=5487;
					out<=51;
				end
				if(in == 3) begin
					state<=3251;
					out<=52;
				end
				if(in == 4) begin
					state<=7140;
					out<=53;
				end
			end
			1598: begin
				if(in == 0) begin
					state<=1599;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=5488;
					out<=56;
				end
				if(in == 3) begin
					state<=3252;
					out<=57;
				end
				if(in == 4) begin
					state<=7141;
					out<=58;
				end
			end
			1599: begin
				if(in == 0) begin
					state<=1600;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=5489;
					out<=61;
				end
				if(in == 3) begin
					state<=3253;
					out<=62;
				end
				if(in == 4) begin
					state<=7142;
					out<=63;
				end
			end
			1600: begin
				if(in == 0) begin
					state<=1601;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=5490;
					out<=66;
				end
				if(in == 3) begin
					state<=3254;
					out<=67;
				end
				if(in == 4) begin
					state<=7143;
					out<=68;
				end
			end
			1601: begin
				if(in == 0) begin
					state<=1602;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=5491;
					out<=71;
				end
				if(in == 3) begin
					state<=3255;
					out<=72;
				end
				if(in == 4) begin
					state<=7144;
					out<=73;
				end
			end
			1602: begin
				if(in == 0) begin
					state<=1603;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=5492;
					out<=76;
				end
				if(in == 3) begin
					state<=3256;
					out<=77;
				end
				if(in == 4) begin
					state<=7145;
					out<=78;
				end
			end
			1603: begin
				if(in == 0) begin
					state<=1604;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=5493;
					out<=81;
				end
				if(in == 3) begin
					state<=3257;
					out<=82;
				end
				if(in == 4) begin
					state<=7146;
					out<=83;
				end
			end
			1604: begin
				if(in == 0) begin
					state<=1605;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=5494;
					out<=86;
				end
				if(in == 3) begin
					state<=3258;
					out<=87;
				end
				if(in == 4) begin
					state<=7147;
					out<=88;
				end
			end
			1605: begin
				if(in == 0) begin
					state<=1606;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=5495;
					out<=91;
				end
				if(in == 3) begin
					state<=3259;
					out<=92;
				end
				if(in == 4) begin
					state<=7148;
					out<=93;
				end
			end
			1606: begin
				if(in == 0) begin
					state<=1607;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=5496;
					out<=96;
				end
				if(in == 3) begin
					state<=3260;
					out<=97;
				end
				if(in == 4) begin
					state<=7149;
					out<=98;
				end
			end
			1607: begin
				if(in == 0) begin
					state<=672;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=4570;
					out<=101;
				end
				if(in == 3) begin
					state<=2670;
					out<=102;
				end
				if(in == 4) begin
					state<=6559;
					out<=103;
				end
			end
			1608: begin
				if(in == 0) begin
					state<=1609;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=5498;
					out<=106;
				end
				if(in == 3) begin
					state<=3510;
					out<=107;
				end
				if(in == 4) begin
					state<=7399;
					out<=108;
				end
			end
			1609: begin
				if(in == 0) begin
					state<=1610;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=5499;
					out<=111;
				end
				if(in == 3) begin
					state<=3511;
					out<=112;
				end
				if(in == 4) begin
					state<=7400;
					out<=113;
				end
			end
			1610: begin
				if(in == 0) begin
					state<=1611;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=5500;
					out<=116;
				end
				if(in == 3) begin
					state<=3512;
					out<=117;
				end
				if(in == 4) begin
					state<=7401;
					out<=118;
				end
			end
			1611: begin
				if(in == 0) begin
					state<=1612;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=5501;
					out<=121;
				end
				if(in == 3) begin
					state<=3513;
					out<=122;
				end
				if(in == 4) begin
					state<=7402;
					out<=123;
				end
			end
			1612: begin
				if(in == 0) begin
					state<=1613;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=5502;
					out<=126;
				end
				if(in == 3) begin
					state<=3514;
					out<=127;
				end
				if(in == 4) begin
					state<=7403;
					out<=128;
				end
			end
			1613: begin
				if(in == 0) begin
					state<=1614;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=5503;
					out<=131;
				end
				if(in == 3) begin
					state<=3515;
					out<=132;
				end
				if(in == 4) begin
					state<=7404;
					out<=133;
				end
			end
			1614: begin
				if(in == 0) begin
					state<=1615;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=5504;
					out<=136;
				end
				if(in == 3) begin
					state<=3516;
					out<=137;
				end
				if(in == 4) begin
					state<=7405;
					out<=138;
				end
			end
			1615: begin
				if(in == 0) begin
					state<=1616;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=5505;
					out<=141;
				end
				if(in == 3) begin
					state<=3517;
					out<=142;
				end
				if(in == 4) begin
					state<=7406;
					out<=143;
				end
			end
			1616: begin
				if(in == 0) begin
					state<=1617;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=5506;
					out<=146;
				end
				if(in == 3) begin
					state<=3518;
					out<=147;
				end
				if(in == 4) begin
					state<=7407;
					out<=148;
				end
			end
			1617: begin
				if(in == 0) begin
					state<=1618;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=5507;
					out<=151;
				end
				if(in == 3) begin
					state<=3519;
					out<=152;
				end
				if(in == 4) begin
					state<=7408;
					out<=153;
				end
			end
			1618: begin
				if(in == 0) begin
					state<=1619;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=5508;
					out<=156;
				end
				if(in == 3) begin
					state<=3520;
					out<=157;
				end
				if(in == 4) begin
					state<=7409;
					out<=158;
				end
			end
			1619: begin
				if(in == 0) begin
					state<=1620;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=5509;
					out<=161;
				end
				if(in == 3) begin
					state<=3521;
					out<=162;
				end
				if(in == 4) begin
					state<=7410;
					out<=163;
				end
			end
			1620: begin
				if(in == 0) begin
					state<=1621;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=5510;
					out<=166;
				end
				if(in == 3) begin
					state<=3522;
					out<=167;
				end
				if(in == 4) begin
					state<=7411;
					out<=168;
				end
			end
			1621: begin
				if(in == 0) begin
					state<=1622;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=5511;
					out<=171;
				end
				if(in == 3) begin
					state<=3523;
					out<=172;
				end
				if(in == 4) begin
					state<=7412;
					out<=173;
				end
			end
			1622: begin
				if(in == 0) begin
					state<=1623;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=5512;
					out<=176;
				end
				if(in == 3) begin
					state<=3524;
					out<=177;
				end
				if(in == 4) begin
					state<=7413;
					out<=178;
				end
			end
			1623: begin
				if(in == 0) begin
					state<=1624;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=5513;
					out<=181;
				end
				if(in == 3) begin
					state<=3525;
					out<=182;
				end
				if(in == 4) begin
					state<=7414;
					out<=183;
				end
			end
			1624: begin
				if(in == 0) begin
					state<=1625;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=5514;
					out<=186;
				end
				if(in == 3) begin
					state<=3526;
					out<=187;
				end
				if(in == 4) begin
					state<=7415;
					out<=188;
				end
			end
			1625: begin
				if(in == 0) begin
					state<=1626;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=5515;
					out<=191;
				end
				if(in == 3) begin
					state<=3527;
					out<=192;
				end
				if(in == 4) begin
					state<=7416;
					out<=193;
				end
			end
			1626: begin
				if(in == 0) begin
					state<=1627;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=5516;
					out<=196;
				end
				if(in == 3) begin
					state<=3528;
					out<=197;
				end
				if(in == 4) begin
					state<=7417;
					out<=198;
				end
			end
			1627: begin
				if(in == 0) begin
					state<=1628;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=5517;
					out<=201;
				end
				if(in == 3) begin
					state<=3529;
					out<=202;
				end
				if(in == 4) begin
					state<=7418;
					out<=203;
				end
			end
			1628: begin
				if(in == 0) begin
					state<=1629;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=5518;
					out<=206;
				end
				if(in == 3) begin
					state<=3530;
					out<=207;
				end
				if(in == 4) begin
					state<=7419;
					out<=208;
				end
			end
			1629: begin
				if(in == 0) begin
					state<=1630;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=5519;
					out<=211;
				end
				if(in == 3) begin
					state<=3531;
					out<=212;
				end
				if(in == 4) begin
					state<=7420;
					out<=213;
				end
			end
			1630: begin
				if(in == 0) begin
					state<=1631;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=5520;
					out<=216;
				end
				if(in == 3) begin
					state<=3532;
					out<=217;
				end
				if(in == 4) begin
					state<=7421;
					out<=218;
				end
			end
			1631: begin
				if(in == 0) begin
					state<=1632;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=5521;
					out<=221;
				end
				if(in == 3) begin
					state<=3533;
					out<=222;
				end
				if(in == 4) begin
					state<=7422;
					out<=223;
				end
			end
			1632: begin
				if(in == 0) begin
					state<=1633;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=5522;
					out<=226;
				end
				if(in == 3) begin
					state<=3534;
					out<=227;
				end
				if(in == 4) begin
					state<=7423;
					out<=228;
				end
			end
			1633: begin
				if(in == 0) begin
					state<=1634;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=5523;
					out<=231;
				end
				if(in == 3) begin
					state<=3535;
					out<=232;
				end
				if(in == 4) begin
					state<=7424;
					out<=233;
				end
			end
			1634: begin
				if(in == 0) begin
					state<=1635;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=5524;
					out<=236;
				end
				if(in == 3) begin
					state<=3536;
					out<=237;
				end
				if(in == 4) begin
					state<=7425;
					out<=238;
				end
			end
			1635: begin
				if(in == 0) begin
					state<=1636;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=5525;
					out<=241;
				end
				if(in == 3) begin
					state<=3537;
					out<=242;
				end
				if(in == 4) begin
					state<=7426;
					out<=243;
				end
			end
			1636: begin
				if(in == 0) begin
					state<=1637;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=5526;
					out<=246;
				end
				if(in == 3) begin
					state<=3538;
					out<=247;
				end
				if(in == 4) begin
					state<=7427;
					out<=248;
				end
			end
			1637: begin
				if(in == 0) begin
					state<=1638;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=5527;
					out<=251;
				end
				if(in == 3) begin
					state<=3539;
					out<=252;
				end
				if(in == 4) begin
					state<=7428;
					out<=253;
				end
			end
			1638: begin
				if(in == 0) begin
					state<=1639;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=5528;
					out<=0;
				end
				if(in == 3) begin
					state<=3540;
					out<=1;
				end
				if(in == 4) begin
					state<=7429;
					out<=2;
				end
			end
			1639: begin
				if(in == 0) begin
					state<=1640;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=5529;
					out<=5;
				end
				if(in == 3) begin
					state<=3541;
					out<=6;
				end
				if(in == 4) begin
					state<=7430;
					out<=7;
				end
			end
			1640: begin
				if(in == 0) begin
					state<=1641;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=5530;
					out<=10;
				end
				if(in == 3) begin
					state<=3542;
					out<=11;
				end
				if(in == 4) begin
					state<=7431;
					out<=12;
				end
			end
			1641: begin
				if(in == 0) begin
					state<=1642;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=5531;
					out<=15;
				end
				if(in == 3) begin
					state<=3543;
					out<=16;
				end
				if(in == 4) begin
					state<=7432;
					out<=17;
				end
			end
			1642: begin
				if(in == 0) begin
					state<=1643;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=5532;
					out<=20;
				end
				if(in == 3) begin
					state<=3544;
					out<=21;
				end
				if(in == 4) begin
					state<=7433;
					out<=22;
				end
			end
			1643: begin
				if(in == 0) begin
					state<=1644;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=5533;
					out<=25;
				end
				if(in == 3) begin
					state<=3545;
					out<=26;
				end
				if(in == 4) begin
					state<=7434;
					out<=27;
				end
			end
			1644: begin
				if(in == 0) begin
					state<=1645;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=5534;
					out<=30;
				end
				if(in == 3) begin
					state<=3546;
					out<=31;
				end
				if(in == 4) begin
					state<=7435;
					out<=32;
				end
			end
			1645: begin
				if(in == 0) begin
					state<=1646;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=5535;
					out<=35;
				end
				if(in == 3) begin
					state<=3547;
					out<=36;
				end
				if(in == 4) begin
					state<=7436;
					out<=37;
				end
			end
			1646: begin
				if(in == 0) begin
					state<=1647;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=5536;
					out<=40;
				end
				if(in == 3) begin
					state<=3548;
					out<=41;
				end
				if(in == 4) begin
					state<=7437;
					out<=42;
				end
			end
			1647: begin
				if(in == 0) begin
					state<=1648;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=5537;
					out<=45;
				end
				if(in == 3) begin
					state<=3549;
					out<=46;
				end
				if(in == 4) begin
					state<=7438;
					out<=47;
				end
			end
			1648: begin
				if(in == 0) begin
					state<=1649;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=5538;
					out<=50;
				end
				if(in == 3) begin
					state<=3550;
					out<=51;
				end
				if(in == 4) begin
					state<=7439;
					out<=52;
				end
			end
			1649: begin
				if(in == 0) begin
					state<=1650;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=5539;
					out<=55;
				end
				if(in == 3) begin
					state<=3551;
					out<=56;
				end
				if(in == 4) begin
					state<=7440;
					out<=57;
				end
			end
			1650: begin
				if(in == 0) begin
					state<=1651;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=5540;
					out<=60;
				end
				if(in == 3) begin
					state<=3552;
					out<=61;
				end
				if(in == 4) begin
					state<=7441;
					out<=62;
				end
			end
			1651: begin
				if(in == 0) begin
					state<=1652;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=5541;
					out<=65;
				end
				if(in == 3) begin
					state<=3553;
					out<=66;
				end
				if(in == 4) begin
					state<=7442;
					out<=67;
				end
			end
			1652: begin
				if(in == 0) begin
					state<=1653;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=5542;
					out<=70;
				end
				if(in == 3) begin
					state<=3554;
					out<=71;
				end
				if(in == 4) begin
					state<=7443;
					out<=72;
				end
			end
			1653: begin
				if(in == 0) begin
					state<=1654;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=5543;
					out<=75;
				end
				if(in == 3) begin
					state<=3555;
					out<=76;
				end
				if(in == 4) begin
					state<=7444;
					out<=77;
				end
			end
			1654: begin
				if(in == 0) begin
					state<=1655;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=5544;
					out<=80;
				end
				if(in == 3) begin
					state<=3556;
					out<=81;
				end
				if(in == 4) begin
					state<=7445;
					out<=82;
				end
			end
			1655: begin
				if(in == 0) begin
					state<=1656;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=5545;
					out<=85;
				end
				if(in == 3) begin
					state<=3557;
					out<=86;
				end
				if(in == 4) begin
					state<=7446;
					out<=87;
				end
			end
			1656: begin
				if(in == 0) begin
					state<=1657;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=5546;
					out<=90;
				end
				if(in == 3) begin
					state<=3558;
					out<=91;
				end
				if(in == 4) begin
					state<=7447;
					out<=92;
				end
			end
			1657: begin
				if(in == 0) begin
					state<=1658;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=5547;
					out<=95;
				end
				if(in == 3) begin
					state<=3559;
					out<=96;
				end
				if(in == 4) begin
					state<=7448;
					out<=97;
				end
			end
			1658: begin
				if(in == 0) begin
					state<=1659;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=5548;
					out<=100;
				end
				if(in == 3) begin
					state<=3560;
					out<=101;
				end
				if(in == 4) begin
					state<=7449;
					out<=102;
				end
			end
			1659: begin
				if(in == 0) begin
					state<=1660;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=5549;
					out<=105;
				end
				if(in == 3) begin
					state<=3561;
					out<=106;
				end
				if(in == 4) begin
					state<=7450;
					out<=107;
				end
			end
			1660: begin
				if(in == 0) begin
					state<=1661;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=5550;
					out<=110;
				end
				if(in == 3) begin
					state<=3562;
					out<=111;
				end
				if(in == 4) begin
					state<=7451;
					out<=112;
				end
			end
			1661: begin
				if(in == 0) begin
					state<=1662;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=5551;
					out<=115;
				end
				if(in == 3) begin
					state<=3563;
					out<=116;
				end
				if(in == 4) begin
					state<=7452;
					out<=117;
				end
			end
			1662: begin
				if(in == 0) begin
					state<=1663;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=5552;
					out<=120;
				end
				if(in == 3) begin
					state<=3564;
					out<=121;
				end
				if(in == 4) begin
					state<=7453;
					out<=122;
				end
			end
			1663: begin
				if(in == 0) begin
					state<=1664;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=5553;
					out<=125;
				end
				if(in == 3) begin
					state<=3565;
					out<=126;
				end
				if(in == 4) begin
					state<=7454;
					out<=127;
				end
			end
			1664: begin
				if(in == 0) begin
					state<=1665;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=5554;
					out<=130;
				end
				if(in == 3) begin
					state<=3566;
					out<=131;
				end
				if(in == 4) begin
					state<=7455;
					out<=132;
				end
			end
			1665: begin
				if(in == 0) begin
					state<=1666;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=5555;
					out<=135;
				end
				if(in == 3) begin
					state<=3567;
					out<=136;
				end
				if(in == 4) begin
					state<=7456;
					out<=137;
				end
			end
			1666: begin
				if(in == 0) begin
					state<=1667;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=5556;
					out<=140;
				end
				if(in == 3) begin
					state<=3568;
					out<=141;
				end
				if(in == 4) begin
					state<=7457;
					out<=142;
				end
			end
			1667: begin
				if(in == 0) begin
					state<=1668;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=5557;
					out<=145;
				end
				if(in == 3) begin
					state<=3569;
					out<=146;
				end
				if(in == 4) begin
					state<=7458;
					out<=147;
				end
			end
			1668: begin
				if(in == 0) begin
					state<=1669;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=5558;
					out<=150;
				end
				if(in == 3) begin
					state<=3570;
					out<=151;
				end
				if(in == 4) begin
					state<=7459;
					out<=152;
				end
			end
			1669: begin
				if(in == 0) begin
					state<=1670;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=5559;
					out<=155;
				end
				if(in == 3) begin
					state<=3571;
					out<=156;
				end
				if(in == 4) begin
					state<=7460;
					out<=157;
				end
			end
			1670: begin
				if(in == 0) begin
					state<=1671;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=5560;
					out<=160;
				end
				if(in == 3) begin
					state<=3572;
					out<=161;
				end
				if(in == 4) begin
					state<=7461;
					out<=162;
				end
			end
			1671: begin
				if(in == 0) begin
					state<=1672;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=5561;
					out<=165;
				end
				if(in == 3) begin
					state<=3573;
					out<=166;
				end
				if(in == 4) begin
					state<=7462;
					out<=167;
				end
			end
			1672: begin
				if(in == 0) begin
					state<=1673;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=5562;
					out<=170;
				end
				if(in == 3) begin
					state<=3574;
					out<=171;
				end
				if(in == 4) begin
					state<=7463;
					out<=172;
				end
			end
			1673: begin
				if(in == 0) begin
					state<=1674;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=5563;
					out<=175;
				end
				if(in == 3) begin
					state<=3575;
					out<=176;
				end
				if(in == 4) begin
					state<=7464;
					out<=177;
				end
			end
			1674: begin
				if(in == 0) begin
					state<=1675;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=5564;
					out<=180;
				end
				if(in == 3) begin
					state<=3576;
					out<=181;
				end
				if(in == 4) begin
					state<=7465;
					out<=182;
				end
			end
			1675: begin
				if(in == 0) begin
					state<=1676;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=5565;
					out<=185;
				end
				if(in == 3) begin
					state<=3577;
					out<=186;
				end
				if(in == 4) begin
					state<=7466;
					out<=187;
				end
			end
			1676: begin
				if(in == 0) begin
					state<=1677;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=5566;
					out<=190;
				end
				if(in == 3) begin
					state<=3578;
					out<=191;
				end
				if(in == 4) begin
					state<=7467;
					out<=192;
				end
			end
			1677: begin
				if(in == 0) begin
					state<=1678;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=5567;
					out<=195;
				end
				if(in == 3) begin
					state<=3579;
					out<=196;
				end
				if(in == 4) begin
					state<=7468;
					out<=197;
				end
			end
			1678: begin
				if(in == 0) begin
					state<=1679;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=5568;
					out<=200;
				end
				if(in == 3) begin
					state<=3580;
					out<=201;
				end
				if(in == 4) begin
					state<=7469;
					out<=202;
				end
			end
			1679: begin
				if(in == 0) begin
					state<=1680;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=5569;
					out<=205;
				end
				if(in == 3) begin
					state<=3581;
					out<=206;
				end
				if(in == 4) begin
					state<=7470;
					out<=207;
				end
			end
			1680: begin
				if(in == 0) begin
					state<=1681;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=5570;
					out<=210;
				end
				if(in == 3) begin
					state<=3582;
					out<=211;
				end
				if(in == 4) begin
					state<=7471;
					out<=212;
				end
			end
			1681: begin
				if(in == 0) begin
					state<=1682;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=5571;
					out<=215;
				end
				if(in == 3) begin
					state<=3583;
					out<=216;
				end
				if(in == 4) begin
					state<=7472;
					out<=217;
				end
			end
			1682: begin
				if(in == 0) begin
					state<=1683;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=5572;
					out<=220;
				end
				if(in == 3) begin
					state<=3584;
					out<=221;
				end
				if(in == 4) begin
					state<=7473;
					out<=222;
				end
			end
			1683: begin
				if(in == 0) begin
					state<=1684;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=5573;
					out<=225;
				end
				if(in == 3) begin
					state<=3585;
					out<=226;
				end
				if(in == 4) begin
					state<=7474;
					out<=227;
				end
			end
			1684: begin
				if(in == 0) begin
					state<=1685;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=5574;
					out<=230;
				end
				if(in == 3) begin
					state<=3586;
					out<=231;
				end
				if(in == 4) begin
					state<=7475;
					out<=232;
				end
			end
			1685: begin
				if(in == 0) begin
					state<=1686;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=5575;
					out<=235;
				end
				if(in == 3) begin
					state<=3587;
					out<=236;
				end
				if(in == 4) begin
					state<=7476;
					out<=237;
				end
			end
			1686: begin
				if(in == 0) begin
					state<=1687;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=5576;
					out<=240;
				end
				if(in == 3) begin
					state<=3588;
					out<=241;
				end
				if(in == 4) begin
					state<=7477;
					out<=242;
				end
			end
			1687: begin
				if(in == 0) begin
					state<=1688;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=5577;
					out<=245;
				end
				if(in == 3) begin
					state<=3589;
					out<=246;
				end
				if(in == 4) begin
					state<=7478;
					out<=247;
				end
			end
			1688: begin
				if(in == 0) begin
					state<=1689;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=5578;
					out<=250;
				end
				if(in == 3) begin
					state<=3590;
					out<=251;
				end
				if(in == 4) begin
					state<=7479;
					out<=252;
				end
			end
			1689: begin
				if(in == 0) begin
					state<=1690;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=5579;
					out<=255;
				end
				if(in == 3) begin
					state<=3591;
					out<=0;
				end
				if(in == 4) begin
					state<=7480;
					out<=1;
				end
			end
			1690: begin
				if(in == 0) begin
					state<=1691;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=5580;
					out<=4;
				end
				if(in == 3) begin
					state<=3592;
					out<=5;
				end
				if(in == 4) begin
					state<=7481;
					out<=6;
				end
			end
			1691: begin
				if(in == 0) begin
					state<=1692;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=5581;
					out<=9;
				end
				if(in == 3) begin
					state<=3593;
					out<=10;
				end
				if(in == 4) begin
					state<=7482;
					out<=11;
				end
			end
			1692: begin
				if(in == 0) begin
					state<=1693;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=5582;
					out<=14;
				end
				if(in == 3) begin
					state<=3594;
					out<=15;
				end
				if(in == 4) begin
					state<=7483;
					out<=16;
				end
			end
			1693: begin
				if(in == 0) begin
					state<=1694;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=5583;
					out<=19;
				end
				if(in == 3) begin
					state<=3595;
					out<=20;
				end
				if(in == 4) begin
					state<=7484;
					out<=21;
				end
			end
			1694: begin
				if(in == 0) begin
					state<=1695;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=5584;
					out<=24;
				end
				if(in == 3) begin
					state<=3596;
					out<=25;
				end
				if(in == 4) begin
					state<=7485;
					out<=26;
				end
			end
			1695: begin
				if(in == 0) begin
					state<=1696;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=5585;
					out<=29;
				end
				if(in == 3) begin
					state<=3597;
					out<=30;
				end
				if(in == 4) begin
					state<=7486;
					out<=31;
				end
			end
			1696: begin
				if(in == 0) begin
					state<=1697;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=5586;
					out<=34;
				end
				if(in == 3) begin
					state<=3598;
					out<=35;
				end
				if(in == 4) begin
					state<=7487;
					out<=36;
				end
			end
			1697: begin
				if(in == 0) begin
					state<=1698;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=5587;
					out<=39;
				end
				if(in == 3) begin
					state<=3599;
					out<=40;
				end
				if(in == 4) begin
					state<=7488;
					out<=41;
				end
			end
			1698: begin
				if(in == 0) begin
					state<=1699;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=5588;
					out<=44;
				end
				if(in == 3) begin
					state<=3600;
					out<=45;
				end
				if(in == 4) begin
					state<=7489;
					out<=46;
				end
			end
			1699: begin
				if(in == 0) begin
					state<=1700;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=5589;
					out<=49;
				end
				if(in == 3) begin
					state<=3601;
					out<=50;
				end
				if(in == 4) begin
					state<=7490;
					out<=51;
				end
			end
			1700: begin
				if(in == 0) begin
					state<=1701;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=5590;
					out<=54;
				end
				if(in == 3) begin
					state<=3602;
					out<=55;
				end
				if(in == 4) begin
					state<=7491;
					out<=56;
				end
			end
			1701: begin
				if(in == 0) begin
					state<=1702;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=5591;
					out<=59;
				end
				if(in == 3) begin
					state<=3603;
					out<=60;
				end
				if(in == 4) begin
					state<=7492;
					out<=61;
				end
			end
			1702: begin
				if(in == 0) begin
					state<=1703;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=5592;
					out<=64;
				end
				if(in == 3) begin
					state<=3604;
					out<=65;
				end
				if(in == 4) begin
					state<=7493;
					out<=66;
				end
			end
			1703: begin
				if(in == 0) begin
					state<=1704;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=5593;
					out<=69;
				end
				if(in == 3) begin
					state<=3605;
					out<=70;
				end
				if(in == 4) begin
					state<=7494;
					out<=71;
				end
			end
			1704: begin
				if(in == 0) begin
					state<=1705;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=5594;
					out<=74;
				end
				if(in == 3) begin
					state<=3606;
					out<=75;
				end
				if(in == 4) begin
					state<=7495;
					out<=76;
				end
			end
			1705: begin
				if(in == 0) begin
					state<=1706;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=5595;
					out<=79;
				end
				if(in == 3) begin
					state<=3607;
					out<=80;
				end
				if(in == 4) begin
					state<=7496;
					out<=81;
				end
			end
			1706: begin
				if(in == 0) begin
					state<=1707;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=5596;
					out<=84;
				end
				if(in == 3) begin
					state<=3608;
					out<=85;
				end
				if(in == 4) begin
					state<=7497;
					out<=86;
				end
			end
			1707: begin
				if(in == 0) begin
					state<=1708;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=5597;
					out<=89;
				end
				if(in == 3) begin
					state<=3609;
					out<=90;
				end
				if(in == 4) begin
					state<=7498;
					out<=91;
				end
			end
			1708: begin
				if(in == 0) begin
					state<=1709;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=5598;
					out<=94;
				end
				if(in == 3) begin
					state<=3610;
					out<=95;
				end
				if(in == 4) begin
					state<=7499;
					out<=96;
				end
			end
			1709: begin
				if(in == 0) begin
					state<=1710;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=5599;
					out<=99;
				end
				if(in == 3) begin
					state<=3611;
					out<=100;
				end
				if(in == 4) begin
					state<=7500;
					out<=101;
				end
			end
			1710: begin
				if(in == 0) begin
					state<=1711;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=5600;
					out<=104;
				end
				if(in == 3) begin
					state<=3612;
					out<=105;
				end
				if(in == 4) begin
					state<=7501;
					out<=106;
				end
			end
			1711: begin
				if(in == 0) begin
					state<=1712;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=5601;
					out<=109;
				end
				if(in == 3) begin
					state<=3613;
					out<=110;
				end
				if(in == 4) begin
					state<=7502;
					out<=111;
				end
			end
			1712: begin
				if(in == 0) begin
					state<=1713;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=5602;
					out<=114;
				end
				if(in == 3) begin
					state<=3614;
					out<=115;
				end
				if(in == 4) begin
					state<=7503;
					out<=116;
				end
			end
			1713: begin
				if(in == 0) begin
					state<=1714;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=5603;
					out<=119;
				end
				if(in == 3) begin
					state<=3615;
					out<=120;
				end
				if(in == 4) begin
					state<=7504;
					out<=121;
				end
			end
			1714: begin
				if(in == 0) begin
					state<=1715;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=5604;
					out<=124;
				end
				if(in == 3) begin
					state<=3616;
					out<=125;
				end
				if(in == 4) begin
					state<=7505;
					out<=126;
				end
			end
			1715: begin
				if(in == 0) begin
					state<=1716;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=5605;
					out<=129;
				end
				if(in == 3) begin
					state<=3617;
					out<=130;
				end
				if(in == 4) begin
					state<=7506;
					out<=131;
				end
			end
			1716: begin
				if(in == 0) begin
					state<=1717;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=5606;
					out<=134;
				end
				if(in == 3) begin
					state<=3618;
					out<=135;
				end
				if(in == 4) begin
					state<=7507;
					out<=136;
				end
			end
			1717: begin
				if(in == 0) begin
					state<=1718;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=5607;
					out<=139;
				end
				if(in == 3) begin
					state<=3619;
					out<=140;
				end
				if(in == 4) begin
					state<=7508;
					out<=141;
				end
			end
			1718: begin
				if(in == 0) begin
					state<=1719;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=5608;
					out<=144;
				end
				if(in == 3) begin
					state<=3620;
					out<=145;
				end
				if(in == 4) begin
					state<=7509;
					out<=146;
				end
			end
			1719: begin
				if(in == 0) begin
					state<=1720;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=5609;
					out<=149;
				end
				if(in == 3) begin
					state<=3621;
					out<=150;
				end
				if(in == 4) begin
					state<=7510;
					out<=151;
				end
			end
			1720: begin
				if(in == 0) begin
					state<=1721;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=5610;
					out<=154;
				end
				if(in == 3) begin
					state<=3622;
					out<=155;
				end
				if(in == 4) begin
					state<=7511;
					out<=156;
				end
			end
			1721: begin
				if(in == 0) begin
					state<=1722;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=5611;
					out<=159;
				end
				if(in == 3) begin
					state<=3623;
					out<=160;
				end
				if(in == 4) begin
					state<=7512;
					out<=161;
				end
			end
			1722: begin
				if(in == 0) begin
					state<=1723;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=5612;
					out<=164;
				end
				if(in == 3) begin
					state<=3624;
					out<=165;
				end
				if(in == 4) begin
					state<=7513;
					out<=166;
				end
			end
			1723: begin
				if(in == 0) begin
					state<=1724;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=5613;
					out<=169;
				end
				if(in == 3) begin
					state<=3625;
					out<=170;
				end
				if(in == 4) begin
					state<=7514;
					out<=171;
				end
			end
			1724: begin
				if(in == 0) begin
					state<=1725;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=5614;
					out<=174;
				end
				if(in == 3) begin
					state<=3626;
					out<=175;
				end
				if(in == 4) begin
					state<=7515;
					out<=176;
				end
			end
			1725: begin
				if(in == 0) begin
					state<=1726;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=5615;
					out<=179;
				end
				if(in == 3) begin
					state<=3627;
					out<=180;
				end
				if(in == 4) begin
					state<=7516;
					out<=181;
				end
			end
			1726: begin
				if(in == 0) begin
					state<=1727;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=5616;
					out<=184;
				end
				if(in == 3) begin
					state<=3628;
					out<=185;
				end
				if(in == 4) begin
					state<=7517;
					out<=186;
				end
			end
			1727: begin
				if(in == 0) begin
					state<=1728;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=5617;
					out<=189;
				end
				if(in == 3) begin
					state<=3629;
					out<=190;
				end
				if(in == 4) begin
					state<=7518;
					out<=191;
				end
			end
			1728: begin
				if(in == 0) begin
					state<=1729;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=5618;
					out<=194;
				end
				if(in == 3) begin
					state<=3630;
					out<=195;
				end
				if(in == 4) begin
					state<=7519;
					out<=196;
				end
			end
			1729: begin
				if(in == 0) begin
					state<=1730;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=5619;
					out<=199;
				end
				if(in == 3) begin
					state<=3631;
					out<=200;
				end
				if(in == 4) begin
					state<=7520;
					out<=201;
				end
			end
			1730: begin
				if(in == 0) begin
					state<=1731;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=5620;
					out<=204;
				end
				if(in == 3) begin
					state<=3632;
					out<=205;
				end
				if(in == 4) begin
					state<=7521;
					out<=206;
				end
			end
			1731: begin
				if(in == 0) begin
					state<=1732;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=5621;
					out<=209;
				end
				if(in == 3) begin
					state<=3633;
					out<=210;
				end
				if(in == 4) begin
					state<=7522;
					out<=211;
				end
			end
			1732: begin
				if(in == 0) begin
					state<=1733;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=5622;
					out<=214;
				end
				if(in == 3) begin
					state<=3634;
					out<=215;
				end
				if(in == 4) begin
					state<=7523;
					out<=216;
				end
			end
			1733: begin
				if(in == 0) begin
					state<=1734;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=5623;
					out<=219;
				end
				if(in == 3) begin
					state<=3635;
					out<=220;
				end
				if(in == 4) begin
					state<=7524;
					out<=221;
				end
			end
			1734: begin
				if(in == 0) begin
					state<=1735;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=5624;
					out<=224;
				end
				if(in == 3) begin
					state<=3636;
					out<=225;
				end
				if(in == 4) begin
					state<=7525;
					out<=226;
				end
			end
			1735: begin
				if(in == 0) begin
					state<=1736;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=5625;
					out<=229;
				end
				if(in == 3) begin
					state<=3637;
					out<=230;
				end
				if(in == 4) begin
					state<=7526;
					out<=231;
				end
			end
			1736: begin
				if(in == 0) begin
					state<=1737;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=5626;
					out<=234;
				end
				if(in == 3) begin
					state<=3638;
					out<=235;
				end
				if(in == 4) begin
					state<=7527;
					out<=236;
				end
			end
			1737: begin
				if(in == 0) begin
					state<=1738;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=5627;
					out<=239;
				end
				if(in == 3) begin
					state<=3639;
					out<=240;
				end
				if(in == 4) begin
					state<=7528;
					out<=241;
				end
			end
			1738: begin
				if(in == 0) begin
					state<=1739;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=5628;
					out<=244;
				end
				if(in == 3) begin
					state<=3640;
					out<=245;
				end
				if(in == 4) begin
					state<=7529;
					out<=246;
				end
			end
			1739: begin
				if(in == 0) begin
					state<=1740;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=5629;
					out<=249;
				end
				if(in == 3) begin
					state<=3641;
					out<=250;
				end
				if(in == 4) begin
					state<=7530;
					out<=251;
				end
			end
			1740: begin
				if(in == 0) begin
					state<=1741;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=5630;
					out<=254;
				end
				if(in == 3) begin
					state<=3642;
					out<=255;
				end
				if(in == 4) begin
					state<=7531;
					out<=0;
				end
			end
			1741: begin
				if(in == 0) begin
					state<=1742;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=5631;
					out<=3;
				end
				if(in == 3) begin
					state<=3643;
					out<=4;
				end
				if(in == 4) begin
					state<=7532;
					out<=5;
				end
			end
			1742: begin
				if(in == 0) begin
					state<=1743;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=5632;
					out<=8;
				end
				if(in == 3) begin
					state<=3644;
					out<=9;
				end
				if(in == 4) begin
					state<=7533;
					out<=10;
				end
			end
			1743: begin
				if(in == 0) begin
					state<=1744;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=5633;
					out<=13;
				end
				if(in == 3) begin
					state<=3645;
					out<=14;
				end
				if(in == 4) begin
					state<=7534;
					out<=15;
				end
			end
			1744: begin
				if(in == 0) begin
					state<=1745;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=5634;
					out<=18;
				end
				if(in == 3) begin
					state<=3646;
					out<=19;
				end
				if(in == 4) begin
					state<=7535;
					out<=20;
				end
			end
			1745: begin
				if(in == 0) begin
					state<=1746;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=5635;
					out<=23;
				end
				if(in == 3) begin
					state<=3647;
					out<=24;
				end
				if(in == 4) begin
					state<=7536;
					out<=25;
				end
			end
			1746: begin
				if(in == 0) begin
					state<=1747;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=5636;
					out<=28;
				end
				if(in == 3) begin
					state<=3648;
					out<=29;
				end
				if(in == 4) begin
					state<=7537;
					out<=30;
				end
			end
			1747: begin
				if(in == 0) begin
					state<=1748;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=5637;
					out<=33;
				end
				if(in == 3) begin
					state<=3649;
					out<=34;
				end
				if(in == 4) begin
					state<=7538;
					out<=35;
				end
			end
			1748: begin
				if(in == 0) begin
					state<=1749;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=5638;
					out<=38;
				end
				if(in == 3) begin
					state<=3650;
					out<=39;
				end
				if(in == 4) begin
					state<=7539;
					out<=40;
				end
			end
			1749: begin
				if(in == 0) begin
					state<=1750;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=5639;
					out<=43;
				end
				if(in == 3) begin
					state<=3651;
					out<=44;
				end
				if(in == 4) begin
					state<=7540;
					out<=45;
				end
			end
			1750: begin
				if(in == 0) begin
					state<=1751;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=5640;
					out<=48;
				end
				if(in == 3) begin
					state<=3652;
					out<=49;
				end
				if(in == 4) begin
					state<=7541;
					out<=50;
				end
			end
			1751: begin
				if(in == 0) begin
					state<=1752;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=5641;
					out<=53;
				end
				if(in == 3) begin
					state<=3653;
					out<=54;
				end
				if(in == 4) begin
					state<=7542;
					out<=55;
				end
			end
			1752: begin
				if(in == 0) begin
					state<=1753;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=5642;
					out<=58;
				end
				if(in == 3) begin
					state<=3654;
					out<=59;
				end
				if(in == 4) begin
					state<=7543;
					out<=60;
				end
			end
			1753: begin
				if(in == 0) begin
					state<=1754;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=5643;
					out<=63;
				end
				if(in == 3) begin
					state<=3655;
					out<=64;
				end
				if(in == 4) begin
					state<=7544;
					out<=65;
				end
			end
			1754: begin
				if(in == 0) begin
					state<=1755;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=5644;
					out<=68;
				end
				if(in == 3) begin
					state<=3656;
					out<=69;
				end
				if(in == 4) begin
					state<=7545;
					out<=70;
				end
			end
			1755: begin
				if(in == 0) begin
					state<=1756;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=5645;
					out<=73;
				end
				if(in == 3) begin
					state<=3657;
					out<=74;
				end
				if(in == 4) begin
					state<=7546;
					out<=75;
				end
			end
			1756: begin
				if(in == 0) begin
					state<=1757;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=5646;
					out<=78;
				end
				if(in == 3) begin
					state<=3658;
					out<=79;
				end
				if(in == 4) begin
					state<=7547;
					out<=80;
				end
			end
			1757: begin
				if(in == 0) begin
					state<=1758;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=5647;
					out<=83;
				end
				if(in == 3) begin
					state<=3659;
					out<=84;
				end
				if(in == 4) begin
					state<=7548;
					out<=85;
				end
			end
			1758: begin
				if(in == 0) begin
					state<=1759;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=5648;
					out<=88;
				end
				if(in == 3) begin
					state<=3660;
					out<=89;
				end
				if(in == 4) begin
					state<=7549;
					out<=90;
				end
			end
			1759: begin
				if(in == 0) begin
					state<=1760;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=5649;
					out<=93;
				end
				if(in == 3) begin
					state<=3661;
					out<=94;
				end
				if(in == 4) begin
					state<=7550;
					out<=95;
				end
			end
			1760: begin
				if(in == 0) begin
					state<=1761;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=5650;
					out<=98;
				end
				if(in == 3) begin
					state<=3662;
					out<=99;
				end
				if(in == 4) begin
					state<=7551;
					out<=100;
				end
			end
			1761: begin
				if(in == 0) begin
					state<=1762;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=5651;
					out<=103;
				end
				if(in == 3) begin
					state<=3663;
					out<=104;
				end
				if(in == 4) begin
					state<=7552;
					out<=105;
				end
			end
			1762: begin
				if(in == 0) begin
					state<=1763;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=5652;
					out<=108;
				end
				if(in == 3) begin
					state<=3664;
					out<=109;
				end
				if(in == 4) begin
					state<=7553;
					out<=110;
				end
			end
			1763: begin
				if(in == 0) begin
					state<=1764;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=5653;
					out<=113;
				end
				if(in == 3) begin
					state<=3665;
					out<=114;
				end
				if(in == 4) begin
					state<=7554;
					out<=115;
				end
			end
			1764: begin
				if(in == 0) begin
					state<=1765;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=5654;
					out<=118;
				end
				if(in == 3) begin
					state<=3666;
					out<=119;
				end
				if(in == 4) begin
					state<=7555;
					out<=120;
				end
			end
			1765: begin
				if(in == 0) begin
					state<=1766;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=5655;
					out<=123;
				end
				if(in == 3) begin
					state<=3667;
					out<=124;
				end
				if(in == 4) begin
					state<=7556;
					out<=125;
				end
			end
			1766: begin
				if(in == 0) begin
					state<=1767;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=5656;
					out<=128;
				end
				if(in == 3) begin
					state<=3668;
					out<=129;
				end
				if(in == 4) begin
					state<=7557;
					out<=130;
				end
			end
			1767: begin
				if(in == 0) begin
					state<=1768;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=5657;
					out<=133;
				end
				if(in == 3) begin
					state<=3669;
					out<=134;
				end
				if(in == 4) begin
					state<=7558;
					out<=135;
				end
			end
			1768: begin
				if(in == 0) begin
					state<=1769;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=5658;
					out<=138;
				end
				if(in == 3) begin
					state<=3670;
					out<=139;
				end
				if(in == 4) begin
					state<=7559;
					out<=140;
				end
			end
			1769: begin
				if(in == 0) begin
					state<=1770;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=5659;
					out<=143;
				end
				if(in == 3) begin
					state<=3671;
					out<=144;
				end
				if(in == 4) begin
					state<=7560;
					out<=145;
				end
			end
			1770: begin
				if(in == 0) begin
					state<=1771;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=5660;
					out<=148;
				end
				if(in == 3) begin
					state<=3672;
					out<=149;
				end
				if(in == 4) begin
					state<=7561;
					out<=150;
				end
			end
			1771: begin
				if(in == 0) begin
					state<=1772;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=5661;
					out<=153;
				end
				if(in == 3) begin
					state<=3673;
					out<=154;
				end
				if(in == 4) begin
					state<=7562;
					out<=155;
				end
			end
			1772: begin
				if(in == 0) begin
					state<=1773;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=5662;
					out<=158;
				end
				if(in == 3) begin
					state<=3674;
					out<=159;
				end
				if(in == 4) begin
					state<=7563;
					out<=160;
				end
			end
			1773: begin
				if(in == 0) begin
					state<=1774;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=5663;
					out<=163;
				end
				if(in == 3) begin
					state<=3675;
					out<=164;
				end
				if(in == 4) begin
					state<=7564;
					out<=165;
				end
			end
			1774: begin
				if(in == 0) begin
					state<=1775;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=5664;
					out<=168;
				end
				if(in == 3) begin
					state<=3676;
					out<=169;
				end
				if(in == 4) begin
					state<=7565;
					out<=170;
				end
			end
			1775: begin
				if(in == 0) begin
					state<=1776;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=5665;
					out<=173;
				end
				if(in == 3) begin
					state<=3677;
					out<=174;
				end
				if(in == 4) begin
					state<=7566;
					out<=175;
				end
			end
			1776: begin
				if(in == 0) begin
					state<=1777;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=5666;
					out<=178;
				end
				if(in == 3) begin
					state<=3678;
					out<=179;
				end
				if(in == 4) begin
					state<=7567;
					out<=180;
				end
			end
			1777: begin
				if(in == 0) begin
					state<=1778;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=5667;
					out<=183;
				end
				if(in == 3) begin
					state<=3679;
					out<=184;
				end
				if(in == 4) begin
					state<=7568;
					out<=185;
				end
			end
			1778: begin
				if(in == 0) begin
					state<=1779;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=5668;
					out<=188;
				end
				if(in == 3) begin
					state<=3680;
					out<=189;
				end
				if(in == 4) begin
					state<=7569;
					out<=190;
				end
			end
			1779: begin
				if(in == 0) begin
					state<=1780;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=5669;
					out<=193;
				end
				if(in == 3) begin
					state<=3681;
					out<=194;
				end
				if(in == 4) begin
					state<=7570;
					out<=195;
				end
			end
			1780: begin
				if(in == 0) begin
					state<=1781;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=5670;
					out<=198;
				end
				if(in == 3) begin
					state<=3682;
					out<=199;
				end
				if(in == 4) begin
					state<=7571;
					out<=200;
				end
			end
			1781: begin
				if(in == 0) begin
					state<=1782;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=5671;
					out<=203;
				end
				if(in == 3) begin
					state<=3683;
					out<=204;
				end
				if(in == 4) begin
					state<=7572;
					out<=205;
				end
			end
			1782: begin
				if(in == 0) begin
					state<=1783;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=5672;
					out<=208;
				end
				if(in == 3) begin
					state<=3684;
					out<=209;
				end
				if(in == 4) begin
					state<=7573;
					out<=210;
				end
			end
			1783: begin
				if(in == 0) begin
					state<=1784;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=5673;
					out<=213;
				end
				if(in == 3) begin
					state<=3685;
					out<=214;
				end
				if(in == 4) begin
					state<=7574;
					out<=215;
				end
			end
			1784: begin
				if(in == 0) begin
					state<=1785;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=5674;
					out<=218;
				end
				if(in == 3) begin
					state<=3686;
					out<=219;
				end
				if(in == 4) begin
					state<=7575;
					out<=220;
				end
			end
			1785: begin
				if(in == 0) begin
					state<=1786;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=5675;
					out<=223;
				end
				if(in == 3) begin
					state<=3687;
					out<=224;
				end
				if(in == 4) begin
					state<=7576;
					out<=225;
				end
			end
			1786: begin
				if(in == 0) begin
					state<=1787;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=5676;
					out<=228;
				end
				if(in == 3) begin
					state<=3688;
					out<=229;
				end
				if(in == 4) begin
					state<=7577;
					out<=230;
				end
			end
			1787: begin
				if(in == 0) begin
					state<=1788;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=5677;
					out<=233;
				end
				if(in == 3) begin
					state<=3689;
					out<=234;
				end
				if(in == 4) begin
					state<=7578;
					out<=235;
				end
			end
			1788: begin
				if(in == 0) begin
					state<=1789;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=5678;
					out<=238;
				end
				if(in == 3) begin
					state<=3690;
					out<=239;
				end
				if(in == 4) begin
					state<=7579;
					out<=240;
				end
			end
			1789: begin
				if(in == 0) begin
					state<=1790;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=5679;
					out<=243;
				end
				if(in == 3) begin
					state<=3691;
					out<=244;
				end
				if(in == 4) begin
					state<=7580;
					out<=245;
				end
			end
			1790: begin
				if(in == 0) begin
					state<=1791;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=5680;
					out<=248;
				end
				if(in == 3) begin
					state<=3692;
					out<=249;
				end
				if(in == 4) begin
					state<=7581;
					out<=250;
				end
			end
			1791: begin
				if(in == 0) begin
					state<=1792;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=5681;
					out<=253;
				end
				if(in == 3) begin
					state<=3693;
					out<=254;
				end
				if(in == 4) begin
					state<=7582;
					out<=255;
				end
			end
			1792: begin
				if(in == 0) begin
					state<=1793;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=5682;
					out<=2;
				end
				if(in == 3) begin
					state<=3694;
					out<=3;
				end
				if(in == 4) begin
					state<=7583;
					out<=4;
				end
			end
			1793: begin
				if(in == 0) begin
					state<=1794;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=5683;
					out<=7;
				end
				if(in == 3) begin
					state<=3695;
					out<=8;
				end
				if(in == 4) begin
					state<=7584;
					out<=9;
				end
			end
			1794: begin
				if(in == 0) begin
					state<=1795;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=5684;
					out<=12;
				end
				if(in == 3) begin
					state<=3696;
					out<=13;
				end
				if(in == 4) begin
					state<=7585;
					out<=14;
				end
			end
			1795: begin
				if(in == 0) begin
					state<=1796;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=5685;
					out<=17;
				end
				if(in == 3) begin
					state<=3697;
					out<=18;
				end
				if(in == 4) begin
					state<=7586;
					out<=19;
				end
			end
			1796: begin
				if(in == 0) begin
					state<=1797;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=5686;
					out<=22;
				end
				if(in == 3) begin
					state<=3698;
					out<=23;
				end
				if(in == 4) begin
					state<=7587;
					out<=24;
				end
			end
			1797: begin
				if(in == 0) begin
					state<=1798;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=5687;
					out<=27;
				end
				if(in == 3) begin
					state<=3699;
					out<=28;
				end
				if(in == 4) begin
					state<=7588;
					out<=29;
				end
			end
			1798: begin
				if(in == 0) begin
					state<=1799;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=5688;
					out<=32;
				end
				if(in == 3) begin
					state<=3700;
					out<=33;
				end
				if(in == 4) begin
					state<=7589;
					out<=34;
				end
			end
			1799: begin
				if(in == 0) begin
					state<=1800;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=5689;
					out<=37;
				end
				if(in == 3) begin
					state<=3701;
					out<=38;
				end
				if(in == 4) begin
					state<=7590;
					out<=39;
				end
			end
			1800: begin
				if(in == 0) begin
					state<=1801;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=5690;
					out<=42;
				end
				if(in == 3) begin
					state<=3702;
					out<=43;
				end
				if(in == 4) begin
					state<=7591;
					out<=44;
				end
			end
			1801: begin
				if(in == 0) begin
					state<=1802;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=5691;
					out<=47;
				end
				if(in == 3) begin
					state<=3703;
					out<=48;
				end
				if(in == 4) begin
					state<=7592;
					out<=49;
				end
			end
			1802: begin
				if(in == 0) begin
					state<=1803;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=5692;
					out<=52;
				end
				if(in == 3) begin
					state<=3704;
					out<=53;
				end
				if(in == 4) begin
					state<=7593;
					out<=54;
				end
			end
			1803: begin
				if(in == 0) begin
					state<=1804;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=5693;
					out<=57;
				end
				if(in == 3) begin
					state<=3705;
					out<=58;
				end
				if(in == 4) begin
					state<=7594;
					out<=59;
				end
			end
			1804: begin
				if(in == 0) begin
					state<=1805;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=5694;
					out<=62;
				end
				if(in == 3) begin
					state<=3706;
					out<=63;
				end
				if(in == 4) begin
					state<=7595;
					out<=64;
				end
			end
			1805: begin
				if(in == 0) begin
					state<=1806;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=5695;
					out<=67;
				end
				if(in == 3) begin
					state<=3707;
					out<=68;
				end
				if(in == 4) begin
					state<=7596;
					out<=69;
				end
			end
			1806: begin
				if(in == 0) begin
					state<=1807;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=5696;
					out<=72;
				end
				if(in == 3) begin
					state<=3708;
					out<=73;
				end
				if(in == 4) begin
					state<=7597;
					out<=74;
				end
			end
			1807: begin
				if(in == 0) begin
					state<=1808;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=5697;
					out<=77;
				end
				if(in == 3) begin
					state<=3709;
					out<=78;
				end
				if(in == 4) begin
					state<=7598;
					out<=79;
				end
			end
			1808: begin
				if(in == 0) begin
					state<=1809;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=5698;
					out<=82;
				end
				if(in == 3) begin
					state<=3710;
					out<=83;
				end
				if(in == 4) begin
					state<=7599;
					out<=84;
				end
			end
			1809: begin
				if(in == 0) begin
					state<=1810;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=5699;
					out<=87;
				end
				if(in == 3) begin
					state<=3711;
					out<=88;
				end
				if(in == 4) begin
					state<=7600;
					out<=89;
				end
			end
			1810: begin
				if(in == 0) begin
					state<=1811;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=5700;
					out<=92;
				end
				if(in == 3) begin
					state<=3712;
					out<=93;
				end
				if(in == 4) begin
					state<=7601;
					out<=94;
				end
			end
			1811: begin
				if(in == 0) begin
					state<=1812;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=5701;
					out<=97;
				end
				if(in == 3) begin
					state<=3713;
					out<=98;
				end
				if(in == 4) begin
					state<=7602;
					out<=99;
				end
			end
			1812: begin
				if(in == 0) begin
					state<=1813;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=5702;
					out<=102;
				end
				if(in == 3) begin
					state<=3714;
					out<=103;
				end
				if(in == 4) begin
					state<=7603;
					out<=104;
				end
			end
			1813: begin
				if(in == 0) begin
					state<=1814;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=5703;
					out<=107;
				end
				if(in == 3) begin
					state<=3715;
					out<=108;
				end
				if(in == 4) begin
					state<=7604;
					out<=109;
				end
			end
			1814: begin
				if(in == 0) begin
					state<=1815;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=5704;
					out<=112;
				end
				if(in == 3) begin
					state<=3716;
					out<=113;
				end
				if(in == 4) begin
					state<=7605;
					out<=114;
				end
			end
			1815: begin
				if(in == 0) begin
					state<=1816;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=5705;
					out<=117;
				end
				if(in == 3) begin
					state<=3717;
					out<=118;
				end
				if(in == 4) begin
					state<=7606;
					out<=119;
				end
			end
			1816: begin
				if(in == 0) begin
					state<=1817;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=5706;
					out<=122;
				end
				if(in == 3) begin
					state<=3718;
					out<=123;
				end
				if(in == 4) begin
					state<=7607;
					out<=124;
				end
			end
			1817: begin
				if(in == 0) begin
					state<=1818;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=5707;
					out<=127;
				end
				if(in == 3) begin
					state<=3719;
					out<=128;
				end
				if(in == 4) begin
					state<=7608;
					out<=129;
				end
			end
			1818: begin
				if(in == 0) begin
					state<=1819;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=5708;
					out<=132;
				end
				if(in == 3) begin
					state<=3720;
					out<=133;
				end
				if(in == 4) begin
					state<=7609;
					out<=134;
				end
			end
			1819: begin
				if(in == 0) begin
					state<=1820;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=5709;
					out<=137;
				end
				if(in == 3) begin
					state<=3721;
					out<=138;
				end
				if(in == 4) begin
					state<=7610;
					out<=139;
				end
			end
			1820: begin
				if(in == 0) begin
					state<=1821;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=5710;
					out<=142;
				end
				if(in == 3) begin
					state<=3722;
					out<=143;
				end
				if(in == 4) begin
					state<=7611;
					out<=144;
				end
			end
			1821: begin
				if(in == 0) begin
					state<=1822;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=5711;
					out<=147;
				end
				if(in == 3) begin
					state<=3723;
					out<=148;
				end
				if(in == 4) begin
					state<=7612;
					out<=149;
				end
			end
			1822: begin
				if(in == 0) begin
					state<=1823;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=5712;
					out<=152;
				end
				if(in == 3) begin
					state<=3724;
					out<=153;
				end
				if(in == 4) begin
					state<=7613;
					out<=154;
				end
			end
			1823: begin
				if(in == 0) begin
					state<=1824;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=5713;
					out<=157;
				end
				if(in == 3) begin
					state<=3725;
					out<=158;
				end
				if(in == 4) begin
					state<=7614;
					out<=159;
				end
			end
			1824: begin
				if(in == 0) begin
					state<=1825;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=5714;
					out<=162;
				end
				if(in == 3) begin
					state<=3726;
					out<=163;
				end
				if(in == 4) begin
					state<=7615;
					out<=164;
				end
			end
			1825: begin
				if(in == 0) begin
					state<=1826;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=5715;
					out<=167;
				end
				if(in == 3) begin
					state<=3727;
					out<=168;
				end
				if(in == 4) begin
					state<=7616;
					out<=169;
				end
			end
			1826: begin
				if(in == 0) begin
					state<=1827;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=5716;
					out<=172;
				end
				if(in == 3) begin
					state<=3728;
					out<=173;
				end
				if(in == 4) begin
					state<=7617;
					out<=174;
				end
			end
			1827: begin
				if(in == 0) begin
					state<=1828;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=5717;
					out<=177;
				end
				if(in == 3) begin
					state<=3729;
					out<=178;
				end
				if(in == 4) begin
					state<=7618;
					out<=179;
				end
			end
			1828: begin
				if(in == 0) begin
					state<=1829;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=5718;
					out<=182;
				end
				if(in == 3) begin
					state<=3730;
					out<=183;
				end
				if(in == 4) begin
					state<=7619;
					out<=184;
				end
			end
			1829: begin
				if(in == 0) begin
					state<=1830;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=5719;
					out<=187;
				end
				if(in == 3) begin
					state<=3731;
					out<=188;
				end
				if(in == 4) begin
					state<=7620;
					out<=189;
				end
			end
			1830: begin
				if(in == 0) begin
					state<=1831;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=5720;
					out<=192;
				end
				if(in == 3) begin
					state<=3732;
					out<=193;
				end
				if(in == 4) begin
					state<=7621;
					out<=194;
				end
			end
			1831: begin
				if(in == 0) begin
					state<=1832;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=5721;
					out<=197;
				end
				if(in == 3) begin
					state<=3733;
					out<=198;
				end
				if(in == 4) begin
					state<=7622;
					out<=199;
				end
			end
			1832: begin
				if(in == 0) begin
					state<=1833;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=5722;
					out<=202;
				end
				if(in == 3) begin
					state<=3734;
					out<=203;
				end
				if(in == 4) begin
					state<=7623;
					out<=204;
				end
			end
			1833: begin
				if(in == 0) begin
					state<=1834;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=5723;
					out<=207;
				end
				if(in == 3) begin
					state<=3735;
					out<=208;
				end
				if(in == 4) begin
					state<=7624;
					out<=209;
				end
			end
			1834: begin
				if(in == 0) begin
					state<=1835;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=5724;
					out<=212;
				end
				if(in == 3) begin
					state<=3736;
					out<=213;
				end
				if(in == 4) begin
					state<=7625;
					out<=214;
				end
			end
			1835: begin
				if(in == 0) begin
					state<=1836;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=5725;
					out<=217;
				end
				if(in == 3) begin
					state<=3737;
					out<=218;
				end
				if(in == 4) begin
					state<=7626;
					out<=219;
				end
			end
			1836: begin
				if(in == 0) begin
					state<=1837;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=5726;
					out<=222;
				end
				if(in == 3) begin
					state<=3738;
					out<=223;
				end
				if(in == 4) begin
					state<=7627;
					out<=224;
				end
			end
			1837: begin
				if(in == 0) begin
					state<=1838;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=5727;
					out<=227;
				end
				if(in == 3) begin
					state<=3739;
					out<=228;
				end
				if(in == 4) begin
					state<=7628;
					out<=229;
				end
			end
			1838: begin
				if(in == 0) begin
					state<=1839;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=5728;
					out<=232;
				end
				if(in == 3) begin
					state<=3740;
					out<=233;
				end
				if(in == 4) begin
					state<=7629;
					out<=234;
				end
			end
			1839: begin
				if(in == 0) begin
					state<=1840;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=5729;
					out<=237;
				end
				if(in == 3) begin
					state<=3741;
					out<=238;
				end
				if(in == 4) begin
					state<=7630;
					out<=239;
				end
			end
			1840: begin
				if(in == 0) begin
					state<=1841;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=5730;
					out<=242;
				end
				if(in == 3) begin
					state<=3742;
					out<=243;
				end
				if(in == 4) begin
					state<=7631;
					out<=244;
				end
			end
			1841: begin
				if(in == 0) begin
					state<=1842;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=5731;
					out<=247;
				end
				if(in == 3) begin
					state<=3743;
					out<=248;
				end
				if(in == 4) begin
					state<=7632;
					out<=249;
				end
			end
			1842: begin
				if(in == 0) begin
					state<=1843;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=5732;
					out<=252;
				end
				if(in == 3) begin
					state<=3744;
					out<=253;
				end
				if(in == 4) begin
					state<=7633;
					out<=254;
				end
			end
			1843: begin
				if(in == 0) begin
					state<=1844;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=5733;
					out<=1;
				end
				if(in == 3) begin
					state<=3745;
					out<=2;
				end
				if(in == 4) begin
					state<=7634;
					out<=3;
				end
			end
			1844: begin
				if(in == 0) begin
					state<=1845;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=5734;
					out<=6;
				end
				if(in == 3) begin
					state<=3746;
					out<=7;
				end
				if(in == 4) begin
					state<=7635;
					out<=8;
				end
			end
			1845: begin
				if(in == 0) begin
					state<=1846;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=5735;
					out<=11;
				end
				if(in == 3) begin
					state<=3747;
					out<=12;
				end
				if(in == 4) begin
					state<=7636;
					out<=13;
				end
			end
			1846: begin
				if(in == 0) begin
					state<=1847;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=5736;
					out<=16;
				end
				if(in == 3) begin
					state<=3748;
					out<=17;
				end
				if(in == 4) begin
					state<=7637;
					out<=18;
				end
			end
			1847: begin
				if(in == 0) begin
					state<=1848;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=5737;
					out<=21;
				end
				if(in == 3) begin
					state<=3749;
					out<=22;
				end
				if(in == 4) begin
					state<=7638;
					out<=23;
				end
			end
			1848: begin
				if(in == 0) begin
					state<=1849;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=5738;
					out<=26;
				end
				if(in == 3) begin
					state<=3750;
					out<=27;
				end
				if(in == 4) begin
					state<=7639;
					out<=28;
				end
			end
			1849: begin
				if(in == 0) begin
					state<=1850;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=5739;
					out<=31;
				end
				if(in == 3) begin
					state<=3751;
					out<=32;
				end
				if(in == 4) begin
					state<=7640;
					out<=33;
				end
			end
			1850: begin
				if(in == 0) begin
					state<=1851;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=5740;
					out<=36;
				end
				if(in == 3) begin
					state<=3752;
					out<=37;
				end
				if(in == 4) begin
					state<=7641;
					out<=38;
				end
			end
			1851: begin
				if(in == 0) begin
					state<=1852;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=5741;
					out<=41;
				end
				if(in == 3) begin
					state<=3753;
					out<=42;
				end
				if(in == 4) begin
					state<=7642;
					out<=43;
				end
			end
			1852: begin
				if(in == 0) begin
					state<=1853;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=5742;
					out<=46;
				end
				if(in == 3) begin
					state<=3754;
					out<=47;
				end
				if(in == 4) begin
					state<=7643;
					out<=48;
				end
			end
			1853: begin
				if(in == 0) begin
					state<=1854;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=5743;
					out<=51;
				end
				if(in == 3) begin
					state<=3755;
					out<=52;
				end
				if(in == 4) begin
					state<=7644;
					out<=53;
				end
			end
			1854: begin
				if(in == 0) begin
					state<=1855;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=5744;
					out<=56;
				end
				if(in == 3) begin
					state<=3756;
					out<=57;
				end
				if(in == 4) begin
					state<=7645;
					out<=58;
				end
			end
			1855: begin
				if(in == 0) begin
					state<=1856;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=5745;
					out<=61;
				end
				if(in == 3) begin
					state<=3757;
					out<=62;
				end
				if(in == 4) begin
					state<=7646;
					out<=63;
				end
			end
			1856: begin
				if(in == 0) begin
					state<=1857;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=5746;
					out<=66;
				end
				if(in == 3) begin
					state<=3758;
					out<=67;
				end
				if(in == 4) begin
					state<=7647;
					out<=68;
				end
			end
			1857: begin
				if(in == 0) begin
					state<=1858;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=5747;
					out<=71;
				end
				if(in == 3) begin
					state<=3759;
					out<=72;
				end
				if(in == 4) begin
					state<=7648;
					out<=73;
				end
			end
			1858: begin
				if(in == 0) begin
					state<=1859;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=5748;
					out<=76;
				end
				if(in == 3) begin
					state<=3760;
					out<=77;
				end
				if(in == 4) begin
					state<=7649;
					out<=78;
				end
			end
			1859: begin
				if(in == 0) begin
					state<=1860;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=5749;
					out<=81;
				end
				if(in == 3) begin
					state<=3761;
					out<=82;
				end
				if(in == 4) begin
					state<=7650;
					out<=83;
				end
			end
			1860: begin
				if(in == 0) begin
					state<=1861;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=5750;
					out<=86;
				end
				if(in == 3) begin
					state<=3762;
					out<=87;
				end
				if(in == 4) begin
					state<=7651;
					out<=88;
				end
			end
			1861: begin
				if(in == 0) begin
					state<=1862;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=5751;
					out<=91;
				end
				if(in == 3) begin
					state<=3763;
					out<=92;
				end
				if(in == 4) begin
					state<=7652;
					out<=93;
				end
			end
			1862: begin
				if(in == 0) begin
					state<=1863;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=5752;
					out<=96;
				end
				if(in == 3) begin
					state<=3764;
					out<=97;
				end
				if(in == 4) begin
					state<=7653;
					out<=98;
				end
			end
			1863: begin
				if(in == 0) begin
					state<=1864;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=5753;
					out<=101;
				end
				if(in == 3) begin
					state<=3765;
					out<=102;
				end
				if(in == 4) begin
					state<=7654;
					out<=103;
				end
			end
			1864: begin
				if(in == 0) begin
					state<=1865;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=5754;
					out<=106;
				end
				if(in == 3) begin
					state<=3766;
					out<=107;
				end
				if(in == 4) begin
					state<=7655;
					out<=108;
				end
			end
			1865: begin
				if(in == 0) begin
					state<=1866;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=5755;
					out<=111;
				end
				if(in == 3) begin
					state<=3767;
					out<=112;
				end
				if(in == 4) begin
					state<=7656;
					out<=113;
				end
			end
			1866: begin
				if(in == 0) begin
					state<=1867;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=5756;
					out<=116;
				end
				if(in == 3) begin
					state<=3768;
					out<=117;
				end
				if(in == 4) begin
					state<=7657;
					out<=118;
				end
			end
			1867: begin
				if(in == 0) begin
					state<=1868;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=5757;
					out<=121;
				end
				if(in == 3) begin
					state<=3769;
					out<=122;
				end
				if(in == 4) begin
					state<=7658;
					out<=123;
				end
			end
			1868: begin
				if(in == 0) begin
					state<=1869;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=5758;
					out<=126;
				end
				if(in == 3) begin
					state<=3770;
					out<=127;
				end
				if(in == 4) begin
					state<=7659;
					out<=128;
				end
			end
			1869: begin
				if(in == 0) begin
					state<=1870;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=5759;
					out<=131;
				end
				if(in == 3) begin
					state<=3771;
					out<=132;
				end
				if(in == 4) begin
					state<=7660;
					out<=133;
				end
			end
			1870: begin
				if(in == 0) begin
					state<=1871;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=5760;
					out<=136;
				end
				if(in == 3) begin
					state<=3772;
					out<=137;
				end
				if(in == 4) begin
					state<=7661;
					out<=138;
				end
			end
			1871: begin
				if(in == 0) begin
					state<=1872;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=5761;
					out<=141;
				end
				if(in == 3) begin
					state<=3773;
					out<=142;
				end
				if(in == 4) begin
					state<=7662;
					out<=143;
				end
			end
			1872: begin
				if(in == 0) begin
					state<=1873;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=5762;
					out<=146;
				end
				if(in == 3) begin
					state<=3774;
					out<=147;
				end
				if(in == 4) begin
					state<=7663;
					out<=148;
				end
			end
			1873: begin
				if(in == 0) begin
					state<=1874;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=5763;
					out<=151;
				end
				if(in == 3) begin
					state<=3775;
					out<=152;
				end
				if(in == 4) begin
					state<=7664;
					out<=153;
				end
			end
			1874: begin
				if(in == 0) begin
					state<=1875;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=5764;
					out<=156;
				end
				if(in == 3) begin
					state<=3776;
					out<=157;
				end
				if(in == 4) begin
					state<=7665;
					out<=158;
				end
			end
			1875: begin
				if(in == 0) begin
					state<=1876;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=5765;
					out<=161;
				end
				if(in == 3) begin
					state<=3777;
					out<=162;
				end
				if(in == 4) begin
					state<=7666;
					out<=163;
				end
			end
			1876: begin
				if(in == 0) begin
					state<=1877;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=5766;
					out<=166;
				end
				if(in == 3) begin
					state<=3778;
					out<=167;
				end
				if(in == 4) begin
					state<=7667;
					out<=168;
				end
			end
			1877: begin
				if(in == 0) begin
					state<=1878;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=5767;
					out<=171;
				end
				if(in == 3) begin
					state<=3779;
					out<=172;
				end
				if(in == 4) begin
					state<=7668;
					out<=173;
				end
			end
			1878: begin
				if(in == 0) begin
					state<=1879;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=5768;
					out<=176;
				end
				if(in == 3) begin
					state<=3780;
					out<=177;
				end
				if(in == 4) begin
					state<=7669;
					out<=178;
				end
			end
			1879: begin
				if(in == 0) begin
					state<=1880;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=5769;
					out<=181;
				end
				if(in == 3) begin
					state<=3781;
					out<=182;
				end
				if(in == 4) begin
					state<=7670;
					out<=183;
				end
			end
			1880: begin
				if(in == 0) begin
					state<=1881;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=5770;
					out<=186;
				end
				if(in == 3) begin
					state<=3782;
					out<=187;
				end
				if(in == 4) begin
					state<=7671;
					out<=188;
				end
			end
			1881: begin
				if(in == 0) begin
					state<=1882;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=5771;
					out<=191;
				end
				if(in == 3) begin
					state<=3783;
					out<=192;
				end
				if(in == 4) begin
					state<=7672;
					out<=193;
				end
			end
			1882: begin
				if(in == 0) begin
					state<=1883;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=5772;
					out<=196;
				end
				if(in == 3) begin
					state<=3784;
					out<=197;
				end
				if(in == 4) begin
					state<=7673;
					out<=198;
				end
			end
			1883: begin
				if(in == 0) begin
					state<=1884;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=5773;
					out<=201;
				end
				if(in == 3) begin
					state<=3785;
					out<=202;
				end
				if(in == 4) begin
					state<=7674;
					out<=203;
				end
			end
			1884: begin
				if(in == 0) begin
					state<=1885;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=5774;
					out<=206;
				end
				if(in == 3) begin
					state<=3786;
					out<=207;
				end
				if(in == 4) begin
					state<=7675;
					out<=208;
				end
			end
			1885: begin
				if(in == 0) begin
					state<=1886;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=5775;
					out<=211;
				end
				if(in == 3) begin
					state<=3787;
					out<=212;
				end
				if(in == 4) begin
					state<=7676;
					out<=213;
				end
			end
			1886: begin
				if(in == 0) begin
					state<=1887;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=5776;
					out<=216;
				end
				if(in == 3) begin
					state<=3788;
					out<=217;
				end
				if(in == 4) begin
					state<=7677;
					out<=218;
				end
			end
			1887: begin
				if(in == 0) begin
					state<=1888;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=5777;
					out<=221;
				end
				if(in == 3) begin
					state<=3789;
					out<=222;
				end
				if(in == 4) begin
					state<=7678;
					out<=223;
				end
			end
			1888: begin
				if(in == 0) begin
					state<=1889;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=5778;
					out<=226;
				end
				if(in == 3) begin
					state<=3790;
					out<=227;
				end
				if(in == 4) begin
					state<=7679;
					out<=228;
				end
			end
			1889: begin
				if(in == 0) begin
					state<=1890;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=5779;
					out<=231;
				end
				if(in == 3) begin
					state<=3791;
					out<=232;
				end
				if(in == 4) begin
					state<=7680;
					out<=233;
				end
			end
			1890: begin
				if(in == 0) begin
					state<=1891;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=5780;
					out<=236;
				end
				if(in == 3) begin
					state<=3792;
					out<=237;
				end
				if(in == 4) begin
					state<=7681;
					out<=238;
				end
			end
			1891: begin
				if(in == 0) begin
					state<=1892;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=5781;
					out<=241;
				end
				if(in == 3) begin
					state<=3793;
					out<=242;
				end
				if(in == 4) begin
					state<=7682;
					out<=243;
				end
			end
			1892: begin
				if(in == 0) begin
					state<=1893;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=5782;
					out<=246;
				end
				if(in == 3) begin
					state<=3794;
					out<=247;
				end
				if(in == 4) begin
					state<=7683;
					out<=248;
				end
			end
			1893: begin
				if(in == 0) begin
					state<=1894;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=5783;
					out<=251;
				end
				if(in == 3) begin
					state<=3795;
					out<=252;
				end
				if(in == 4) begin
					state<=7684;
					out<=253;
				end
			end
			1894: begin
				if(in == 0) begin
					state<=1895;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=5784;
					out<=0;
				end
				if(in == 3) begin
					state<=3796;
					out<=1;
				end
				if(in == 4) begin
					state<=7685;
					out<=2;
				end
			end
			1895: begin
				if(in == 0) begin
					state<=1896;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=5785;
					out<=5;
				end
				if(in == 3) begin
					state<=3797;
					out<=6;
				end
				if(in == 4) begin
					state<=7686;
					out<=7;
				end
			end
			1896: begin
				if(in == 0) begin
					state<=1897;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=5786;
					out<=10;
				end
				if(in == 3) begin
					state<=3798;
					out<=11;
				end
				if(in == 4) begin
					state<=7687;
					out<=12;
				end
			end
			1897: begin
				if(in == 0) begin
					state<=1898;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=5787;
					out<=15;
				end
				if(in == 3) begin
					state<=3799;
					out<=16;
				end
				if(in == 4) begin
					state<=7688;
					out<=17;
				end
			end
			1898: begin
				if(in == 0) begin
					state<=1899;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=5788;
					out<=20;
				end
				if(in == 3) begin
					state<=3800;
					out<=21;
				end
				if(in == 4) begin
					state<=7689;
					out<=22;
				end
			end
			1899: begin
				if(in == 0) begin
					state<=1900;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=5789;
					out<=25;
				end
				if(in == 3) begin
					state<=3801;
					out<=26;
				end
				if(in == 4) begin
					state<=7690;
					out<=27;
				end
			end
			1900: begin
				if(in == 0) begin
					state<=1901;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=5790;
					out<=30;
				end
				if(in == 3) begin
					state<=3802;
					out<=31;
				end
				if(in == 4) begin
					state<=7691;
					out<=32;
				end
			end
			1901: begin
				if(in == 0) begin
					state<=1902;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=5791;
					out<=35;
				end
				if(in == 3) begin
					state<=3803;
					out<=36;
				end
				if(in == 4) begin
					state<=7692;
					out<=37;
				end
			end
			1902: begin
				if(in == 0) begin
					state<=1903;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=5792;
					out<=40;
				end
				if(in == 3) begin
					state<=3804;
					out<=41;
				end
				if(in == 4) begin
					state<=7693;
					out<=42;
				end
			end
			1903: begin
				if(in == 0) begin
					state<=1904;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=5793;
					out<=45;
				end
				if(in == 3) begin
					state<=3805;
					out<=46;
				end
				if(in == 4) begin
					state<=7694;
					out<=47;
				end
			end
			1904: begin
				if(in == 0) begin
					state<=1905;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=5794;
					out<=50;
				end
				if(in == 3) begin
					state<=3806;
					out<=51;
				end
				if(in == 4) begin
					state<=7695;
					out<=52;
				end
			end
			1905: begin
				if(in == 0) begin
					state<=1906;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=5795;
					out<=55;
				end
				if(in == 3) begin
					state<=3807;
					out<=56;
				end
				if(in == 4) begin
					state<=7696;
					out<=57;
				end
			end
			1906: begin
				if(in == 0) begin
					state<=1907;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=5796;
					out<=60;
				end
				if(in == 3) begin
					state<=3808;
					out<=61;
				end
				if(in == 4) begin
					state<=7697;
					out<=62;
				end
			end
			1907: begin
				if(in == 0) begin
					state<=1908;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=5797;
					out<=65;
				end
				if(in == 3) begin
					state<=3809;
					out<=66;
				end
				if(in == 4) begin
					state<=7698;
					out<=67;
				end
			end
			1908: begin
				if(in == 0) begin
					state<=1909;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=5798;
					out<=70;
				end
				if(in == 3) begin
					state<=3810;
					out<=71;
				end
				if(in == 4) begin
					state<=7699;
					out<=72;
				end
			end
			1909: begin
				if(in == 0) begin
					state<=1910;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=5799;
					out<=75;
				end
				if(in == 3) begin
					state<=3811;
					out<=76;
				end
				if(in == 4) begin
					state<=7700;
					out<=77;
				end
			end
			1910: begin
				if(in == 0) begin
					state<=1911;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=5800;
					out<=80;
				end
				if(in == 3) begin
					state<=3812;
					out<=81;
				end
				if(in == 4) begin
					state<=7701;
					out<=82;
				end
			end
			1911: begin
				if(in == 0) begin
					state<=1912;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=5801;
					out<=85;
				end
				if(in == 3) begin
					state<=3813;
					out<=86;
				end
				if(in == 4) begin
					state<=7702;
					out<=87;
				end
			end
			1912: begin
				if(in == 0) begin
					state<=1913;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=5802;
					out<=90;
				end
				if(in == 3) begin
					state<=3814;
					out<=91;
				end
				if(in == 4) begin
					state<=7703;
					out<=92;
				end
			end
			1913: begin
				if(in == 0) begin
					state<=1914;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=5803;
					out<=95;
				end
				if(in == 3) begin
					state<=3815;
					out<=96;
				end
				if(in == 4) begin
					state<=7704;
					out<=97;
				end
			end
			1914: begin
				if(in == 0) begin
					state<=1915;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=5804;
					out<=100;
				end
				if(in == 3) begin
					state<=3816;
					out<=101;
				end
				if(in == 4) begin
					state<=7705;
					out<=102;
				end
			end
			1915: begin
				if(in == 0) begin
					state<=1916;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=5805;
					out<=105;
				end
				if(in == 3) begin
					state<=3817;
					out<=106;
				end
				if(in == 4) begin
					state<=7706;
					out<=107;
				end
			end
			1916: begin
				if(in == 0) begin
					state<=1917;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=5806;
					out<=110;
				end
				if(in == 3) begin
					state<=3818;
					out<=111;
				end
				if(in == 4) begin
					state<=7707;
					out<=112;
				end
			end
			1917: begin
				if(in == 0) begin
					state<=1918;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=5807;
					out<=115;
				end
				if(in == 3) begin
					state<=3819;
					out<=116;
				end
				if(in == 4) begin
					state<=7708;
					out<=117;
				end
			end
			1918: begin
				if(in == 0) begin
					state<=1919;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=5808;
					out<=120;
				end
				if(in == 3) begin
					state<=3820;
					out<=121;
				end
				if(in == 4) begin
					state<=7709;
					out<=122;
				end
			end
			1919: begin
				if(in == 0) begin
					state<=1920;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=5809;
					out<=125;
				end
				if(in == 3) begin
					state<=3821;
					out<=126;
				end
				if(in == 4) begin
					state<=7710;
					out<=127;
				end
			end
			1920: begin
				if(in == 0) begin
					state<=1921;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=5810;
					out<=130;
				end
				if(in == 3) begin
					state<=3822;
					out<=131;
				end
				if(in == 4) begin
					state<=7711;
					out<=132;
				end
			end
			1921: begin
				if(in == 0) begin
					state<=1922;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=5811;
					out<=135;
				end
				if(in == 3) begin
					state<=3823;
					out<=136;
				end
				if(in == 4) begin
					state<=7712;
					out<=137;
				end
			end
			1922: begin
				if(in == 0) begin
					state<=1923;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=5812;
					out<=140;
				end
				if(in == 3) begin
					state<=3824;
					out<=141;
				end
				if(in == 4) begin
					state<=7713;
					out<=142;
				end
			end
			1923: begin
				if(in == 0) begin
					state<=1924;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=5813;
					out<=145;
				end
				if(in == 3) begin
					state<=3825;
					out<=146;
				end
				if(in == 4) begin
					state<=7714;
					out<=147;
				end
			end
			1924: begin
				if(in == 0) begin
					state<=1925;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=5814;
					out<=150;
				end
				if(in == 3) begin
					state<=3826;
					out<=151;
				end
				if(in == 4) begin
					state<=7715;
					out<=152;
				end
			end
			1925: begin
				if(in == 0) begin
					state<=1926;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=5815;
					out<=155;
				end
				if(in == 3) begin
					state<=3827;
					out<=156;
				end
				if(in == 4) begin
					state<=7716;
					out<=157;
				end
			end
			1926: begin
				if(in == 0) begin
					state<=1927;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=5816;
					out<=160;
				end
				if(in == 3) begin
					state<=3828;
					out<=161;
				end
				if(in == 4) begin
					state<=7717;
					out<=162;
				end
			end
			1927: begin
				if(in == 0) begin
					state<=1928;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=5817;
					out<=165;
				end
				if(in == 3) begin
					state<=3829;
					out<=166;
				end
				if(in == 4) begin
					state<=7718;
					out<=167;
				end
			end
			1928: begin
				if(in == 0) begin
					state<=1929;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=5818;
					out<=170;
				end
				if(in == 3) begin
					state<=3830;
					out<=171;
				end
				if(in == 4) begin
					state<=7719;
					out<=172;
				end
			end
			1929: begin
				if(in == 0) begin
					state<=1930;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=5819;
					out<=175;
				end
				if(in == 3) begin
					state<=3831;
					out<=176;
				end
				if(in == 4) begin
					state<=7720;
					out<=177;
				end
			end
			1930: begin
				if(in == 0) begin
					state<=1931;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=5820;
					out<=180;
				end
				if(in == 3) begin
					state<=3832;
					out<=181;
				end
				if(in == 4) begin
					state<=7721;
					out<=182;
				end
			end
			1931: begin
				if(in == 0) begin
					state<=1932;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=5821;
					out<=185;
				end
				if(in == 3) begin
					state<=3833;
					out<=186;
				end
				if(in == 4) begin
					state<=7722;
					out<=187;
				end
			end
			1932: begin
				if(in == 0) begin
					state<=1933;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=5822;
					out<=190;
				end
				if(in == 3) begin
					state<=3834;
					out<=191;
				end
				if(in == 4) begin
					state<=7723;
					out<=192;
				end
			end
			1933: begin
				if(in == 0) begin
					state<=1934;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=5823;
					out<=195;
				end
				if(in == 3) begin
					state<=3835;
					out<=196;
				end
				if(in == 4) begin
					state<=7724;
					out<=197;
				end
			end
			1934: begin
				if(in == 0) begin
					state<=1935;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=5824;
					out<=200;
				end
				if(in == 3) begin
					state<=3836;
					out<=201;
				end
				if(in == 4) begin
					state<=7725;
					out<=202;
				end
			end
			1935: begin
				if(in == 0) begin
					state<=1936;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=5825;
					out<=205;
				end
				if(in == 3) begin
					state<=3837;
					out<=206;
				end
				if(in == 4) begin
					state<=7726;
					out<=207;
				end
			end
			1936: begin
				if(in == 0) begin
					state<=1937;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=5826;
					out<=210;
				end
				if(in == 3) begin
					state<=3838;
					out<=211;
				end
				if(in == 4) begin
					state<=7727;
					out<=212;
				end
			end
			1937: begin
				if(in == 0) begin
					state<=1938;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=5827;
					out<=215;
				end
				if(in == 3) begin
					state<=3839;
					out<=216;
				end
				if(in == 4) begin
					state<=7728;
					out<=217;
				end
			end
			1938: begin
				if(in == 0) begin
					state<=1939;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=5828;
					out<=220;
				end
				if(in == 3) begin
					state<=3840;
					out<=221;
				end
				if(in == 4) begin
					state<=7729;
					out<=222;
				end
			end
			1939: begin
				if(in == 0) begin
					state<=1940;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=5829;
					out<=225;
				end
				if(in == 3) begin
					state<=3841;
					out<=226;
				end
				if(in == 4) begin
					state<=7730;
					out<=227;
				end
			end
			1940: begin
				if(in == 0) begin
					state<=1941;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=5830;
					out<=230;
				end
				if(in == 3) begin
					state<=3842;
					out<=231;
				end
				if(in == 4) begin
					state<=7731;
					out<=232;
				end
			end
			1941: begin
				if(in == 0) begin
					state<=1942;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=5831;
					out<=235;
				end
				if(in == 3) begin
					state<=3843;
					out<=236;
				end
				if(in == 4) begin
					state<=7732;
					out<=237;
				end
			end
			1942: begin
				if(in == 0) begin
					state<=1943;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=5832;
					out<=240;
				end
				if(in == 3) begin
					state<=3844;
					out<=241;
				end
				if(in == 4) begin
					state<=7733;
					out<=242;
				end
			end
			1943: begin
				if(in == 0) begin
					state<=1944;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=5833;
					out<=245;
				end
				if(in == 3) begin
					state<=3845;
					out<=246;
				end
				if(in == 4) begin
					state<=7734;
					out<=247;
				end
			end
			1944: begin
				if(in == 0) begin
					state<=1945;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=5834;
					out<=250;
				end
				if(in == 3) begin
					state<=3846;
					out<=251;
				end
				if(in == 4) begin
					state<=7735;
					out<=252;
				end
			end
			1945: begin
				if(in == 0) begin
					state<=1946;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=5835;
					out<=255;
				end
				if(in == 3) begin
					state<=3847;
					out<=0;
				end
				if(in == 4) begin
					state<=7736;
					out<=1;
				end
			end
			1946: begin
				if(in == 0) begin
					state<=1947;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=5836;
					out<=4;
				end
				if(in == 3) begin
					state<=3848;
					out<=5;
				end
				if(in == 4) begin
					state<=7737;
					out<=6;
				end
			end
			1947: begin
				if(in == 0) begin
					state<=1948;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=5837;
					out<=9;
				end
				if(in == 3) begin
					state<=3849;
					out<=10;
				end
				if(in == 4) begin
					state<=7738;
					out<=11;
				end
			end
			1948: begin
				if(in == 0) begin
					state<=1949;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=5838;
					out<=14;
				end
				if(in == 3) begin
					state<=3850;
					out<=15;
				end
				if(in == 4) begin
					state<=7739;
					out<=16;
				end
			end
			1949: begin
				if(in == 0) begin
					state<=1950;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=5839;
					out<=19;
				end
				if(in == 3) begin
					state<=3851;
					out<=20;
				end
				if(in == 4) begin
					state<=7740;
					out<=21;
				end
			end
			1950: begin
				if(in == 0) begin
					state<=1951;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=5840;
					out<=24;
				end
				if(in == 3) begin
					state<=3852;
					out<=25;
				end
				if(in == 4) begin
					state<=7741;
					out<=26;
				end
			end
			1951: begin
				if(in == 0) begin
					state<=1952;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=5841;
					out<=29;
				end
				if(in == 3) begin
					state<=3853;
					out<=30;
				end
				if(in == 4) begin
					state<=7742;
					out<=31;
				end
			end
			1952: begin
				if(in == 0) begin
					state<=1953;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=5842;
					out<=34;
				end
				if(in == 3) begin
					state<=3854;
					out<=35;
				end
				if(in == 4) begin
					state<=7743;
					out<=36;
				end
			end
			1953: begin
				if(in == 0) begin
					state<=1954;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=5843;
					out<=39;
				end
				if(in == 3) begin
					state<=3855;
					out<=40;
				end
				if(in == 4) begin
					state<=7744;
					out<=41;
				end
			end
			1954: begin
				if(in == 0) begin
					state<=1955;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=5844;
					out<=44;
				end
				if(in == 3) begin
					state<=3856;
					out<=45;
				end
				if(in == 4) begin
					state<=7745;
					out<=46;
				end
			end
			1955: begin
				if(in == 0) begin
					state<=1956;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=5845;
					out<=49;
				end
				if(in == 3) begin
					state<=3857;
					out<=50;
				end
				if(in == 4) begin
					state<=7746;
					out<=51;
				end
			end
			1956: begin
				if(in == 0) begin
					state<=1957;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=5846;
					out<=54;
				end
				if(in == 3) begin
					state<=3858;
					out<=55;
				end
				if(in == 4) begin
					state<=7747;
					out<=56;
				end
			end
			1957: begin
				if(in == 0) begin
					state<=1958;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=5847;
					out<=59;
				end
				if(in == 3) begin
					state<=3859;
					out<=60;
				end
				if(in == 4) begin
					state<=7748;
					out<=61;
				end
			end
			1958: begin
				if(in == 0) begin
					state<=1959;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=5848;
					out<=64;
				end
				if(in == 3) begin
					state<=3860;
					out<=65;
				end
				if(in == 4) begin
					state<=7749;
					out<=66;
				end
			end
			1959: begin
				if(in == 0) begin
					state<=1960;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=5849;
					out<=69;
				end
				if(in == 3) begin
					state<=3861;
					out<=70;
				end
				if(in == 4) begin
					state<=7750;
					out<=71;
				end
			end
			1960: begin
				if(in == 0) begin
					state<=1961;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=5850;
					out<=74;
				end
				if(in == 3) begin
					state<=3862;
					out<=75;
				end
				if(in == 4) begin
					state<=7751;
					out<=76;
				end
			end
			1961: begin
				if(in == 0) begin
					state<=1962;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=5851;
					out<=79;
				end
				if(in == 3) begin
					state<=3863;
					out<=80;
				end
				if(in == 4) begin
					state<=7752;
					out<=81;
				end
			end
			1962: begin
				if(in == 0) begin
					state<=1963;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=5852;
					out<=84;
				end
				if(in == 3) begin
					state<=3864;
					out<=85;
				end
				if(in == 4) begin
					state<=7753;
					out<=86;
				end
			end
			1963: begin
				if(in == 0) begin
					state<=1964;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=5853;
					out<=89;
				end
				if(in == 3) begin
					state<=3865;
					out<=90;
				end
				if(in == 4) begin
					state<=7754;
					out<=91;
				end
			end
			1964: begin
				if(in == 0) begin
					state<=1965;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=5854;
					out<=94;
				end
				if(in == 3) begin
					state<=3866;
					out<=95;
				end
				if(in == 4) begin
					state<=7755;
					out<=96;
				end
			end
			1965: begin
				if(in == 0) begin
					state<=1966;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=5855;
					out<=99;
				end
				if(in == 3) begin
					state<=3867;
					out<=100;
				end
				if(in == 4) begin
					state<=7756;
					out<=101;
				end
			end
			1966: begin
				if(in == 0) begin
					state<=1967;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=5856;
					out<=104;
				end
				if(in == 3) begin
					state<=3868;
					out<=105;
				end
				if(in == 4) begin
					state<=7757;
					out<=106;
				end
			end
			1967: begin
				if(in == 0) begin
					state<=1968;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=5857;
					out<=109;
				end
				if(in == 3) begin
					state<=3869;
					out<=110;
				end
				if(in == 4) begin
					state<=7758;
					out<=111;
				end
			end
			1968: begin
				if(in == 0) begin
					state<=1969;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=5858;
					out<=114;
				end
				if(in == 3) begin
					state<=3870;
					out<=115;
				end
				if(in == 4) begin
					state<=7759;
					out<=116;
				end
			end
			1969: begin
				if(in == 0) begin
					state<=1970;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=5859;
					out<=119;
				end
				if(in == 3) begin
					state<=3871;
					out<=120;
				end
				if(in == 4) begin
					state<=7760;
					out<=121;
				end
			end
			1970: begin
				if(in == 0) begin
					state<=1971;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=5860;
					out<=124;
				end
				if(in == 3) begin
					state<=3872;
					out<=125;
				end
				if(in == 4) begin
					state<=7761;
					out<=126;
				end
			end
			1971: begin
				if(in == 0) begin
					state<=1972;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=5861;
					out<=129;
				end
				if(in == 3) begin
					state<=3873;
					out<=130;
				end
				if(in == 4) begin
					state<=7762;
					out<=131;
				end
			end
			1972: begin
				if(in == 0) begin
					state<=1973;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=5862;
					out<=134;
				end
				if(in == 3) begin
					state<=3874;
					out<=135;
				end
				if(in == 4) begin
					state<=7763;
					out<=136;
				end
			end
			1973: begin
				if(in == 0) begin
					state<=1974;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=5863;
					out<=139;
				end
				if(in == 3) begin
					state<=3875;
					out<=140;
				end
				if(in == 4) begin
					state<=7764;
					out<=141;
				end
			end
			1974: begin
				if(in == 0) begin
					state<=1975;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=5864;
					out<=144;
				end
				if(in == 3) begin
					state<=3876;
					out<=145;
				end
				if(in == 4) begin
					state<=7765;
					out<=146;
				end
			end
			1975: begin
				if(in == 0) begin
					state<=1976;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=5865;
					out<=149;
				end
				if(in == 3) begin
					state<=3877;
					out<=150;
				end
				if(in == 4) begin
					state<=7766;
					out<=151;
				end
			end
			1976: begin
				if(in == 0) begin
					state<=1977;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=5866;
					out<=154;
				end
				if(in == 3) begin
					state<=3878;
					out<=155;
				end
				if(in == 4) begin
					state<=7767;
					out<=156;
				end
			end
			1977: begin
				if(in == 0) begin
					state<=1978;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=5867;
					out<=159;
				end
				if(in == 3) begin
					state<=3879;
					out<=160;
				end
				if(in == 4) begin
					state<=7768;
					out<=161;
				end
			end
			1978: begin
				if(in == 0) begin
					state<=1979;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=5868;
					out<=164;
				end
				if(in == 3) begin
					state<=3880;
					out<=165;
				end
				if(in == 4) begin
					state<=7769;
					out<=166;
				end
			end
			1979: begin
				if(in == 0) begin
					state<=1980;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=5869;
					out<=169;
				end
				if(in == 3) begin
					state<=3881;
					out<=170;
				end
				if(in == 4) begin
					state<=7770;
					out<=171;
				end
			end
			1980: begin
				if(in == 0) begin
					state<=1981;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=5870;
					out<=174;
				end
				if(in == 3) begin
					state<=3882;
					out<=175;
				end
				if(in == 4) begin
					state<=7771;
					out<=176;
				end
			end
			1981: begin
				if(in == 0) begin
					state<=1982;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=5871;
					out<=179;
				end
				if(in == 3) begin
					state<=3883;
					out<=180;
				end
				if(in == 4) begin
					state<=7772;
					out<=181;
				end
			end
			1982: begin
				if(in == 0) begin
					state<=1983;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=5872;
					out<=184;
				end
				if(in == 3) begin
					state<=3884;
					out<=185;
				end
				if(in == 4) begin
					state<=7773;
					out<=186;
				end
			end
			1983: begin
				if(in == 0) begin
					state<=1984;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=5873;
					out<=189;
				end
				if(in == 3) begin
					state<=3885;
					out<=190;
				end
				if(in == 4) begin
					state<=7774;
					out<=191;
				end
			end
			1984: begin
				if(in == 0) begin
					state<=1985;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=5874;
					out<=194;
				end
				if(in == 3) begin
					state<=3886;
					out<=195;
				end
				if(in == 4) begin
					state<=7775;
					out<=196;
				end
			end
			1985: begin
				if(in == 0) begin
					state<=1986;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=5875;
					out<=199;
				end
				if(in == 3) begin
					state<=3887;
					out<=200;
				end
				if(in == 4) begin
					state<=7776;
					out<=201;
				end
			end
			1986: begin
				if(in == 0) begin
					state<=1987;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=5876;
					out<=204;
				end
				if(in == 3) begin
					state<=3888;
					out<=205;
				end
				if(in == 4) begin
					state<=7777;
					out<=206;
				end
			end
			1987: begin
				if(in == 0) begin
					state<=1988;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=5877;
					out<=209;
				end
				if(in == 3) begin
					state<=3889;
					out<=210;
				end
				if(in == 4) begin
					state<=7778;
					out<=211;
				end
			end
			1988: begin
				if(in == 0) begin
					state<=1989;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=5878;
					out<=214;
				end
				if(in == 3) begin
					state<=3890;
					out<=215;
				end
				if(in == 4) begin
					state<=7779;
					out<=216;
				end
			end
			1989: begin
				if(in == 0) begin
					state<=1990;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=5879;
					out<=219;
				end
				if(in == 3) begin
					state<=3891;
					out<=220;
				end
				if(in == 4) begin
					state<=7780;
					out<=221;
				end
			end
			1990: begin
				if(in == 0) begin
					state<=1991;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=5880;
					out<=224;
				end
				if(in == 3) begin
					state<=3892;
					out<=225;
				end
				if(in == 4) begin
					state<=7781;
					out<=226;
				end
			end
			1991: begin
				if(in == 0) begin
					state<=1992;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=5881;
					out<=229;
				end
				if(in == 3) begin
					state<=3893;
					out<=230;
				end
				if(in == 4) begin
					state<=7782;
					out<=231;
				end
			end
			1992: begin
				if(in == 0) begin
					state<=1993;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=5882;
					out<=234;
				end
				if(in == 3) begin
					state<=3894;
					out<=235;
				end
				if(in == 4) begin
					state<=7783;
					out<=236;
				end
			end
			1993: begin
				if(in == 0) begin
					state<=1994;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=5883;
					out<=239;
				end
				if(in == 3) begin
					state<=3895;
					out<=240;
				end
				if(in == 4) begin
					state<=7784;
					out<=241;
				end
			end
			1994: begin
				if(in == 0) begin
					state<=1995;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=5884;
					out<=244;
				end
				if(in == 3) begin
					state<=3896;
					out<=245;
				end
				if(in == 4) begin
					state<=7785;
					out<=246;
				end
			end
			1995: begin
				if(in == 0) begin
					state<=1996;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=5885;
					out<=249;
				end
				if(in == 3) begin
					state<=3897;
					out<=250;
				end
				if(in == 4) begin
					state<=7786;
					out<=251;
				end
			end
			1996: begin
				if(in == 0) begin
					state<=1997;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=5886;
					out<=254;
				end
				if(in == 3) begin
					state<=3898;
					out<=255;
				end
				if(in == 4) begin
					state<=7787;
					out<=0;
				end
			end
			1997: begin
				if(in == 0) begin
					state<=1998;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=5887;
					out<=3;
				end
				if(in == 3) begin
					state<=2275;
					out<=4;
				end
				if(in == 4) begin
					state<=6164;
					out<=5;
				end
			end
			1998: begin
				if(in == 0) begin
					state<=900;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=4798;
					out<=8;
				end
				if(in == 3) begin
					state<=2276;
					out<=9;
				end
				if(in == 4) begin
					state<=6165;
					out<=10;
				end
			end
			1999: begin
				if(in == 0) begin
					state<=2000;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=5889;
					out<=13;
				end
				if(in == 3) begin
					state<=2;
					out<=14;
				end
				if(in == 4) begin
					state<=3900;
					out<=15;
				end
			end
			2000: begin
				if(in == 0) begin
					state<=2001;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=5890;
					out<=18;
				end
				if(in == 3) begin
					state<=3;
					out<=19;
				end
				if(in == 4) begin
					state<=3901;
					out<=20;
				end
			end
			2001: begin
				if(in == 0) begin
					state<=2002;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=5891;
					out<=23;
				end
				if(in == 3) begin
					state<=4;
					out<=24;
				end
				if(in == 4) begin
					state<=3902;
					out<=25;
				end
			end
			2002: begin
				if(in == 0) begin
					state<=2003;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=5892;
					out<=28;
				end
				if(in == 3) begin
					state<=5;
					out<=29;
				end
				if(in == 4) begin
					state<=3903;
					out<=30;
				end
			end
			2003: begin
				if(in == 0) begin
					state<=2004;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=5893;
					out<=33;
				end
				if(in == 3) begin
					state<=6;
					out<=34;
				end
				if(in == 4) begin
					state<=3904;
					out<=35;
				end
			end
			2004: begin
				if(in == 0) begin
					state<=2005;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=5894;
					out<=38;
				end
				if(in == 3) begin
					state<=7;
					out<=39;
				end
				if(in == 4) begin
					state<=3905;
					out<=40;
				end
			end
			2005: begin
				if(in == 0) begin
					state<=2006;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=5895;
					out<=43;
				end
				if(in == 3) begin
					state<=8;
					out<=44;
				end
				if(in == 4) begin
					state<=3906;
					out<=45;
				end
			end
			2006: begin
				if(in == 0) begin
					state<=2007;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=5896;
					out<=48;
				end
				if(in == 3) begin
					state<=9;
					out<=49;
				end
				if(in == 4) begin
					state<=3907;
					out<=50;
				end
			end
			2007: begin
				if(in == 0) begin
					state<=2008;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=5897;
					out<=53;
				end
				if(in == 3) begin
					state<=10;
					out<=54;
				end
				if(in == 4) begin
					state<=3908;
					out<=55;
				end
			end
			2008: begin
				if(in == 0) begin
					state<=2009;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=5898;
					out<=58;
				end
				if(in == 3) begin
					state<=11;
					out<=59;
				end
				if(in == 4) begin
					state<=3909;
					out<=60;
				end
			end
			2009: begin
				if(in == 0) begin
					state<=2010;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=5899;
					out<=63;
				end
				if(in == 3) begin
					state<=12;
					out<=64;
				end
				if(in == 4) begin
					state<=3910;
					out<=65;
				end
			end
			2010: begin
				if(in == 0) begin
					state<=2011;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=5900;
					out<=68;
				end
				if(in == 3) begin
					state<=13;
					out<=69;
				end
				if(in == 4) begin
					state<=3911;
					out<=70;
				end
			end
			2011: begin
				if(in == 0) begin
					state<=2012;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=5901;
					out<=73;
				end
				if(in == 3) begin
					state<=14;
					out<=74;
				end
				if(in == 4) begin
					state<=3912;
					out<=75;
				end
			end
			2012: begin
				if(in == 0) begin
					state<=2013;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=5902;
					out<=78;
				end
				if(in == 3) begin
					state<=15;
					out<=79;
				end
				if(in == 4) begin
					state<=3913;
					out<=80;
				end
			end
			2013: begin
				if(in == 0) begin
					state<=2014;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=5903;
					out<=83;
				end
				if(in == 3) begin
					state<=16;
					out<=84;
				end
				if(in == 4) begin
					state<=3914;
					out<=85;
				end
			end
			2014: begin
				if(in == 0) begin
					state<=2015;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=5904;
					out<=88;
				end
				if(in == 3) begin
					state<=17;
					out<=89;
				end
				if(in == 4) begin
					state<=3915;
					out<=90;
				end
			end
			2015: begin
				if(in == 0) begin
					state<=2016;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=5905;
					out<=93;
				end
				if(in == 3) begin
					state<=18;
					out<=94;
				end
				if(in == 4) begin
					state<=3916;
					out<=95;
				end
			end
			2016: begin
				if(in == 0) begin
					state<=2017;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=5906;
					out<=98;
				end
				if(in == 3) begin
					state<=19;
					out<=99;
				end
				if(in == 4) begin
					state<=3917;
					out<=100;
				end
			end
			2017: begin
				if(in == 0) begin
					state<=2018;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=5907;
					out<=103;
				end
				if(in == 3) begin
					state<=20;
					out<=104;
				end
				if(in == 4) begin
					state<=3918;
					out<=105;
				end
			end
			2018: begin
				if(in == 0) begin
					state<=2019;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=5908;
					out<=108;
				end
				if(in == 3) begin
					state<=21;
					out<=109;
				end
				if(in == 4) begin
					state<=3919;
					out<=110;
				end
			end
			2019: begin
				if(in == 0) begin
					state<=2020;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=5909;
					out<=113;
				end
				if(in == 3) begin
					state<=22;
					out<=114;
				end
				if(in == 4) begin
					state<=3920;
					out<=115;
				end
			end
			2020: begin
				if(in == 0) begin
					state<=2021;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=5910;
					out<=118;
				end
				if(in == 3) begin
					state<=23;
					out<=119;
				end
				if(in == 4) begin
					state<=3921;
					out<=120;
				end
			end
			2021: begin
				if(in == 0) begin
					state<=2022;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=5911;
					out<=123;
				end
				if(in == 3) begin
					state<=24;
					out<=124;
				end
				if(in == 4) begin
					state<=3922;
					out<=125;
				end
			end
			2022: begin
				if(in == 0) begin
					state<=2023;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=5912;
					out<=128;
				end
				if(in == 3) begin
					state<=25;
					out<=129;
				end
				if(in == 4) begin
					state<=3923;
					out<=130;
				end
			end
			2023: begin
				if(in == 0) begin
					state<=2024;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=5913;
					out<=133;
				end
				if(in == 3) begin
					state<=26;
					out<=134;
				end
				if(in == 4) begin
					state<=3924;
					out<=135;
				end
			end
			2024: begin
				if(in == 0) begin
					state<=2025;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=5914;
					out<=138;
				end
				if(in == 3) begin
					state<=27;
					out<=139;
				end
				if(in == 4) begin
					state<=3925;
					out<=140;
				end
			end
			2025: begin
				if(in == 0) begin
					state<=2026;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=5915;
					out<=143;
				end
				if(in == 3) begin
					state<=28;
					out<=144;
				end
				if(in == 4) begin
					state<=3926;
					out<=145;
				end
			end
			2026: begin
				if(in == 0) begin
					state<=2027;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=5916;
					out<=148;
				end
				if(in == 3) begin
					state<=29;
					out<=149;
				end
				if(in == 4) begin
					state<=3927;
					out<=150;
				end
			end
			2027: begin
				if(in == 0) begin
					state<=2028;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=5917;
					out<=153;
				end
				if(in == 3) begin
					state<=30;
					out<=154;
				end
				if(in == 4) begin
					state<=3928;
					out<=155;
				end
			end
			2028: begin
				if(in == 0) begin
					state<=2029;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=5918;
					out<=158;
				end
				if(in == 3) begin
					state<=31;
					out<=159;
				end
				if(in == 4) begin
					state<=3929;
					out<=160;
				end
			end
			2029: begin
				if(in == 0) begin
					state<=2030;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=5919;
					out<=163;
				end
				if(in == 3) begin
					state<=32;
					out<=164;
				end
				if(in == 4) begin
					state<=3930;
					out<=165;
				end
			end
			2030: begin
				if(in == 0) begin
					state<=2031;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=5920;
					out<=168;
				end
				if(in == 3) begin
					state<=33;
					out<=169;
				end
				if(in == 4) begin
					state<=3931;
					out<=170;
				end
			end
			2031: begin
				if(in == 0) begin
					state<=2032;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=5921;
					out<=173;
				end
				if(in == 3) begin
					state<=34;
					out<=174;
				end
				if(in == 4) begin
					state<=3932;
					out<=175;
				end
			end
			2032: begin
				if(in == 0) begin
					state<=2033;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=5922;
					out<=178;
				end
				if(in == 3) begin
					state<=35;
					out<=179;
				end
				if(in == 4) begin
					state<=3933;
					out<=180;
				end
			end
			2033: begin
				if(in == 0) begin
					state<=2034;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=5923;
					out<=183;
				end
				if(in == 3) begin
					state<=36;
					out<=184;
				end
				if(in == 4) begin
					state<=3934;
					out<=185;
				end
			end
			2034: begin
				if(in == 0) begin
					state<=2035;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=5924;
					out<=188;
				end
				if(in == 3) begin
					state<=37;
					out<=189;
				end
				if(in == 4) begin
					state<=3935;
					out<=190;
				end
			end
			2035: begin
				if(in == 0) begin
					state<=2036;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=5925;
					out<=193;
				end
				if(in == 3) begin
					state<=38;
					out<=194;
				end
				if(in == 4) begin
					state<=3936;
					out<=195;
				end
			end
			2036: begin
				if(in == 0) begin
					state<=2037;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=5926;
					out<=198;
				end
				if(in == 3) begin
					state<=39;
					out<=199;
				end
				if(in == 4) begin
					state<=3937;
					out<=200;
				end
			end
			2037: begin
				if(in == 0) begin
					state<=2038;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=5927;
					out<=203;
				end
				if(in == 3) begin
					state<=40;
					out<=204;
				end
				if(in == 4) begin
					state<=3938;
					out<=205;
				end
			end
			2038: begin
				if(in == 0) begin
					state<=2039;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=5928;
					out<=208;
				end
				if(in == 3) begin
					state<=41;
					out<=209;
				end
				if(in == 4) begin
					state<=3939;
					out<=210;
				end
			end
			2039: begin
				if(in == 0) begin
					state<=2040;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=5929;
					out<=213;
				end
				if(in == 3) begin
					state<=42;
					out<=214;
				end
				if(in == 4) begin
					state<=3940;
					out<=215;
				end
			end
			2040: begin
				if(in == 0) begin
					state<=2041;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=5930;
					out<=218;
				end
				if(in == 3) begin
					state<=43;
					out<=219;
				end
				if(in == 4) begin
					state<=3941;
					out<=220;
				end
			end
			2041: begin
				if(in == 0) begin
					state<=2042;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=5931;
					out<=223;
				end
				if(in == 3) begin
					state<=44;
					out<=224;
				end
				if(in == 4) begin
					state<=3942;
					out<=225;
				end
			end
			2042: begin
				if(in == 0) begin
					state<=2043;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=5932;
					out<=228;
				end
				if(in == 3) begin
					state<=45;
					out<=229;
				end
				if(in == 4) begin
					state<=3943;
					out<=230;
				end
			end
			2043: begin
				if(in == 0) begin
					state<=2044;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=5933;
					out<=233;
				end
				if(in == 3) begin
					state<=46;
					out<=234;
				end
				if(in == 4) begin
					state<=3944;
					out<=235;
				end
			end
			2044: begin
				if(in == 0) begin
					state<=2045;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=5934;
					out<=238;
				end
				if(in == 3) begin
					state<=47;
					out<=239;
				end
				if(in == 4) begin
					state<=3945;
					out<=240;
				end
			end
			2045: begin
				if(in == 0) begin
					state<=2046;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=5935;
					out<=243;
				end
				if(in == 3) begin
					state<=48;
					out<=244;
				end
				if(in == 4) begin
					state<=3946;
					out<=245;
				end
			end
			2046: begin
				if(in == 0) begin
					state<=2047;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=5936;
					out<=248;
				end
				if(in == 3) begin
					state<=49;
					out<=249;
				end
				if(in == 4) begin
					state<=3947;
					out<=250;
				end
			end
			2047: begin
				if(in == 0) begin
					state<=2048;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=5937;
					out<=253;
				end
				if(in == 3) begin
					state<=50;
					out<=254;
				end
				if(in == 4) begin
					state<=3948;
					out<=255;
				end
			end
			2048: begin
				if(in == 0) begin
					state<=3261;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=7150;
					out<=2;
				end
				if(in == 3) begin
					state<=1329;
					out<=3;
				end
				if(in == 4) begin
					state<=5218;
					out<=4;
				end
			end
			2049: begin
				if(in == 0) begin
					state<=2050;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=5939;
					out<=7;
				end
				if(in == 3) begin
					state<=52;
					out<=8;
				end
				if(in == 4) begin
					state<=3950;
					out<=9;
				end
			end
			2050: begin
				if(in == 0) begin
					state<=2051;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=5940;
					out<=12;
				end
				if(in == 3) begin
					state<=53;
					out<=13;
				end
				if(in == 4) begin
					state<=3951;
					out<=14;
				end
			end
			2051: begin
				if(in == 0) begin
					state<=2052;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=5941;
					out<=17;
				end
				if(in == 3) begin
					state<=54;
					out<=18;
				end
				if(in == 4) begin
					state<=3952;
					out<=19;
				end
			end
			2052: begin
				if(in == 0) begin
					state<=2053;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=5942;
					out<=22;
				end
				if(in == 3) begin
					state<=55;
					out<=23;
				end
				if(in == 4) begin
					state<=3953;
					out<=24;
				end
			end
			2053: begin
				if(in == 0) begin
					state<=2054;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=5943;
					out<=27;
				end
				if(in == 3) begin
					state<=56;
					out<=28;
				end
				if(in == 4) begin
					state<=3954;
					out<=29;
				end
			end
			2054: begin
				if(in == 0) begin
					state<=2055;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=5944;
					out<=32;
				end
				if(in == 3) begin
					state<=57;
					out<=33;
				end
				if(in == 4) begin
					state<=3955;
					out<=34;
				end
			end
			2055: begin
				if(in == 0) begin
					state<=2056;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=5945;
					out<=37;
				end
				if(in == 3) begin
					state<=58;
					out<=38;
				end
				if(in == 4) begin
					state<=3956;
					out<=39;
				end
			end
			2056: begin
				if(in == 0) begin
					state<=2057;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=5946;
					out<=42;
				end
				if(in == 3) begin
					state<=59;
					out<=43;
				end
				if(in == 4) begin
					state<=3957;
					out<=44;
				end
			end
			2057: begin
				if(in == 0) begin
					state<=2058;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=5947;
					out<=47;
				end
				if(in == 3) begin
					state<=60;
					out<=48;
				end
				if(in == 4) begin
					state<=3958;
					out<=49;
				end
			end
			2058: begin
				if(in == 0) begin
					state<=2059;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=5948;
					out<=52;
				end
				if(in == 3) begin
					state<=61;
					out<=53;
				end
				if(in == 4) begin
					state<=3959;
					out<=54;
				end
			end
			2059: begin
				if(in == 0) begin
					state<=2060;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=5949;
					out<=57;
				end
				if(in == 3) begin
					state<=62;
					out<=58;
				end
				if(in == 4) begin
					state<=3960;
					out<=59;
				end
			end
			2060: begin
				if(in == 0) begin
					state<=2061;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=5950;
					out<=62;
				end
				if(in == 3) begin
					state<=63;
					out<=63;
				end
				if(in == 4) begin
					state<=3961;
					out<=64;
				end
			end
			2061: begin
				if(in == 0) begin
					state<=2062;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=5951;
					out<=67;
				end
				if(in == 3) begin
					state<=64;
					out<=68;
				end
				if(in == 4) begin
					state<=3962;
					out<=69;
				end
			end
			2062: begin
				if(in == 0) begin
					state<=2063;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=5952;
					out<=72;
				end
				if(in == 3) begin
					state<=65;
					out<=73;
				end
				if(in == 4) begin
					state<=3963;
					out<=74;
				end
			end
			2063: begin
				if(in == 0) begin
					state<=2064;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=5953;
					out<=77;
				end
				if(in == 3) begin
					state<=66;
					out<=78;
				end
				if(in == 4) begin
					state<=3964;
					out<=79;
				end
			end
			2064: begin
				if(in == 0) begin
					state<=2065;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=5954;
					out<=82;
				end
				if(in == 3) begin
					state<=67;
					out<=83;
				end
				if(in == 4) begin
					state<=3965;
					out<=84;
				end
			end
			2065: begin
				if(in == 0) begin
					state<=2066;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=5955;
					out<=87;
				end
				if(in == 3) begin
					state<=68;
					out<=88;
				end
				if(in == 4) begin
					state<=3966;
					out<=89;
				end
			end
			2066: begin
				if(in == 0) begin
					state<=2067;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=5956;
					out<=92;
				end
				if(in == 3) begin
					state<=69;
					out<=93;
				end
				if(in == 4) begin
					state<=3967;
					out<=94;
				end
			end
			2067: begin
				if(in == 0) begin
					state<=2068;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=5957;
					out<=97;
				end
				if(in == 3) begin
					state<=70;
					out<=98;
				end
				if(in == 4) begin
					state<=3968;
					out<=99;
				end
			end
			2068: begin
				if(in == 0) begin
					state<=2069;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=5958;
					out<=102;
				end
				if(in == 3) begin
					state<=71;
					out<=103;
				end
				if(in == 4) begin
					state<=3969;
					out<=104;
				end
			end
			2069: begin
				if(in == 0) begin
					state<=2070;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=5959;
					out<=107;
				end
				if(in == 3) begin
					state<=72;
					out<=108;
				end
				if(in == 4) begin
					state<=3970;
					out<=109;
				end
			end
			2070: begin
				if(in == 0) begin
					state<=2071;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=5960;
					out<=112;
				end
				if(in == 3) begin
					state<=73;
					out<=113;
				end
				if(in == 4) begin
					state<=3971;
					out<=114;
				end
			end
			2071: begin
				if(in == 0) begin
					state<=2072;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=5961;
					out<=117;
				end
				if(in == 3) begin
					state<=74;
					out<=118;
				end
				if(in == 4) begin
					state<=3972;
					out<=119;
				end
			end
			2072: begin
				if(in == 0) begin
					state<=2073;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=5962;
					out<=122;
				end
				if(in == 3) begin
					state<=75;
					out<=123;
				end
				if(in == 4) begin
					state<=3973;
					out<=124;
				end
			end
			2073: begin
				if(in == 0) begin
					state<=2074;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=5963;
					out<=127;
				end
				if(in == 3) begin
					state<=76;
					out<=128;
				end
				if(in == 4) begin
					state<=3974;
					out<=129;
				end
			end
			2074: begin
				if(in == 0) begin
					state<=2075;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=5964;
					out<=132;
				end
				if(in == 3) begin
					state<=77;
					out<=133;
				end
				if(in == 4) begin
					state<=3975;
					out<=134;
				end
			end
			2075: begin
				if(in == 0) begin
					state<=2076;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=5965;
					out<=137;
				end
				if(in == 3) begin
					state<=78;
					out<=138;
				end
				if(in == 4) begin
					state<=3976;
					out<=139;
				end
			end
			2076: begin
				if(in == 0) begin
					state<=2077;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=5966;
					out<=142;
				end
				if(in == 3) begin
					state<=79;
					out<=143;
				end
				if(in == 4) begin
					state<=3977;
					out<=144;
				end
			end
			2077: begin
				if(in == 0) begin
					state<=2078;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=5967;
					out<=147;
				end
				if(in == 3) begin
					state<=80;
					out<=148;
				end
				if(in == 4) begin
					state<=3978;
					out<=149;
				end
			end
			2078: begin
				if(in == 0) begin
					state<=2079;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=5968;
					out<=152;
				end
				if(in == 3) begin
					state<=81;
					out<=153;
				end
				if(in == 4) begin
					state<=3979;
					out<=154;
				end
			end
			2079: begin
				if(in == 0) begin
					state<=2080;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=5969;
					out<=157;
				end
				if(in == 3) begin
					state<=82;
					out<=158;
				end
				if(in == 4) begin
					state<=3980;
					out<=159;
				end
			end
			2080: begin
				if(in == 0) begin
					state<=2081;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=5970;
					out<=162;
				end
				if(in == 3) begin
					state<=83;
					out<=163;
				end
				if(in == 4) begin
					state<=3981;
					out<=164;
				end
			end
			2081: begin
				if(in == 0) begin
					state<=2082;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=5971;
					out<=167;
				end
				if(in == 3) begin
					state<=84;
					out<=168;
				end
				if(in == 4) begin
					state<=3982;
					out<=169;
				end
			end
			2082: begin
				if(in == 0) begin
					state<=2083;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=5972;
					out<=172;
				end
				if(in == 3) begin
					state<=85;
					out<=173;
				end
				if(in == 4) begin
					state<=3983;
					out<=174;
				end
			end
			2083: begin
				if(in == 0) begin
					state<=2084;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=5973;
					out<=177;
				end
				if(in == 3) begin
					state<=86;
					out<=178;
				end
				if(in == 4) begin
					state<=3984;
					out<=179;
				end
			end
			2084: begin
				if(in == 0) begin
					state<=2085;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=5974;
					out<=182;
				end
				if(in == 3) begin
					state<=87;
					out<=183;
				end
				if(in == 4) begin
					state<=3985;
					out<=184;
				end
			end
			2085: begin
				if(in == 0) begin
					state<=2086;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=5975;
					out<=187;
				end
				if(in == 3) begin
					state<=88;
					out<=188;
				end
				if(in == 4) begin
					state<=3986;
					out<=189;
				end
			end
			2086: begin
				if(in == 0) begin
					state<=2087;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=5976;
					out<=192;
				end
				if(in == 3) begin
					state<=89;
					out<=193;
				end
				if(in == 4) begin
					state<=3987;
					out<=194;
				end
			end
			2087: begin
				if(in == 0) begin
					state<=2088;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=5977;
					out<=197;
				end
				if(in == 3) begin
					state<=90;
					out<=198;
				end
				if(in == 4) begin
					state<=3988;
					out<=199;
				end
			end
			2088: begin
				if(in == 0) begin
					state<=2089;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=5978;
					out<=202;
				end
				if(in == 3) begin
					state<=91;
					out<=203;
				end
				if(in == 4) begin
					state<=3989;
					out<=204;
				end
			end
			2089: begin
				if(in == 0) begin
					state<=2090;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=5979;
					out<=207;
				end
				if(in == 3) begin
					state<=92;
					out<=208;
				end
				if(in == 4) begin
					state<=3990;
					out<=209;
				end
			end
			2090: begin
				if(in == 0) begin
					state<=2091;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=5980;
					out<=212;
				end
				if(in == 3) begin
					state<=93;
					out<=213;
				end
				if(in == 4) begin
					state<=3991;
					out<=214;
				end
			end
			2091: begin
				if(in == 0) begin
					state<=2092;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=5981;
					out<=217;
				end
				if(in == 3) begin
					state<=94;
					out<=218;
				end
				if(in == 4) begin
					state<=3992;
					out<=219;
				end
			end
			2092: begin
				if(in == 0) begin
					state<=2093;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=5982;
					out<=222;
				end
				if(in == 3) begin
					state<=95;
					out<=223;
				end
				if(in == 4) begin
					state<=3993;
					out<=224;
				end
			end
			2093: begin
				if(in == 0) begin
					state<=2094;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=5983;
					out<=227;
				end
				if(in == 3) begin
					state<=96;
					out<=228;
				end
				if(in == 4) begin
					state<=3994;
					out<=229;
				end
			end
			2094: begin
				if(in == 0) begin
					state<=2095;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=5984;
					out<=232;
				end
				if(in == 3) begin
					state<=97;
					out<=233;
				end
				if(in == 4) begin
					state<=3995;
					out<=234;
				end
			end
			2095: begin
				if(in == 0) begin
					state<=2096;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=5985;
					out<=237;
				end
				if(in == 3) begin
					state<=98;
					out<=238;
				end
				if(in == 4) begin
					state<=3996;
					out<=239;
				end
			end
			2096: begin
				if(in == 0) begin
					state<=2097;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=5986;
					out<=242;
				end
				if(in == 3) begin
					state<=99;
					out<=243;
				end
				if(in == 4) begin
					state<=3997;
					out<=244;
				end
			end
			2097: begin
				if(in == 0) begin
					state<=2098;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=5987;
					out<=247;
				end
				if(in == 3) begin
					state<=100;
					out<=248;
				end
				if(in == 4) begin
					state<=3998;
					out<=249;
				end
			end
			2098: begin
				if(in == 0) begin
					state<=2099;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=5988;
					out<=252;
				end
				if(in == 3) begin
					state<=101;
					out<=253;
				end
				if(in == 4) begin
					state<=3999;
					out<=254;
				end
			end
			2099: begin
				if(in == 0) begin
					state<=2100;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=5989;
					out<=1;
				end
				if(in == 3) begin
					state<=102;
					out<=2;
				end
				if(in == 4) begin
					state<=4000;
					out<=3;
				end
			end
			2100: begin
				if(in == 0) begin
					state<=2101;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=5990;
					out<=6;
				end
				if(in == 3) begin
					state<=103;
					out<=7;
				end
				if(in == 4) begin
					state<=4001;
					out<=8;
				end
			end
			2101: begin
				if(in == 0) begin
					state<=2102;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=5991;
					out<=11;
				end
				if(in == 3) begin
					state<=104;
					out<=12;
				end
				if(in == 4) begin
					state<=4002;
					out<=13;
				end
			end
			2102: begin
				if(in == 0) begin
					state<=2103;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=5992;
					out<=16;
				end
				if(in == 3) begin
					state<=105;
					out<=17;
				end
				if(in == 4) begin
					state<=4003;
					out<=18;
				end
			end
			2103: begin
				if(in == 0) begin
					state<=2104;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=5993;
					out<=21;
				end
				if(in == 3) begin
					state<=106;
					out<=22;
				end
				if(in == 4) begin
					state<=4004;
					out<=23;
				end
			end
			2104: begin
				if(in == 0) begin
					state<=2105;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=5994;
					out<=26;
				end
				if(in == 3) begin
					state<=107;
					out<=27;
				end
				if(in == 4) begin
					state<=4005;
					out<=28;
				end
			end
			2105: begin
				if(in == 0) begin
					state<=2106;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=5995;
					out<=31;
				end
				if(in == 3) begin
					state<=108;
					out<=32;
				end
				if(in == 4) begin
					state<=4006;
					out<=33;
				end
			end
			2106: begin
				if(in == 0) begin
					state<=2107;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=5996;
					out<=36;
				end
				if(in == 3) begin
					state<=109;
					out<=37;
				end
				if(in == 4) begin
					state<=4007;
					out<=38;
				end
			end
			2107: begin
				if(in == 0) begin
					state<=2108;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=5997;
					out<=41;
				end
				if(in == 3) begin
					state<=110;
					out<=42;
				end
				if(in == 4) begin
					state<=4008;
					out<=43;
				end
			end
			2108: begin
				if(in == 0) begin
					state<=2109;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=5998;
					out<=46;
				end
				if(in == 3) begin
					state<=111;
					out<=47;
				end
				if(in == 4) begin
					state<=4009;
					out<=48;
				end
			end
			2109: begin
				if(in == 0) begin
					state<=2110;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=5999;
					out<=51;
				end
				if(in == 3) begin
					state<=112;
					out<=52;
				end
				if(in == 4) begin
					state<=4010;
					out<=53;
				end
			end
			2110: begin
				if(in == 0) begin
					state<=2111;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=6000;
					out<=56;
				end
				if(in == 3) begin
					state<=113;
					out<=57;
				end
				if(in == 4) begin
					state<=4011;
					out<=58;
				end
			end
			2111: begin
				if(in == 0) begin
					state<=2112;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=6001;
					out<=61;
				end
				if(in == 3) begin
					state<=114;
					out<=62;
				end
				if(in == 4) begin
					state<=4012;
					out<=63;
				end
			end
			2112: begin
				if(in == 0) begin
					state<=2113;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=6002;
					out<=66;
				end
				if(in == 3) begin
					state<=115;
					out<=67;
				end
				if(in == 4) begin
					state<=4013;
					out<=68;
				end
			end
			2113: begin
				if(in == 0) begin
					state<=2114;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=6003;
					out<=71;
				end
				if(in == 3) begin
					state<=116;
					out<=72;
				end
				if(in == 4) begin
					state<=4014;
					out<=73;
				end
			end
			2114: begin
				if(in == 0) begin
					state<=2115;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=6004;
					out<=76;
				end
				if(in == 3) begin
					state<=117;
					out<=77;
				end
				if(in == 4) begin
					state<=4015;
					out<=78;
				end
			end
			2115: begin
				if(in == 0) begin
					state<=2116;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=6005;
					out<=81;
				end
				if(in == 3) begin
					state<=118;
					out<=82;
				end
				if(in == 4) begin
					state<=4016;
					out<=83;
				end
			end
			2116: begin
				if(in == 0) begin
					state<=2117;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=6006;
					out<=86;
				end
				if(in == 3) begin
					state<=119;
					out<=87;
				end
				if(in == 4) begin
					state<=4017;
					out<=88;
				end
			end
			2117: begin
				if(in == 0) begin
					state<=3292;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=7181;
					out<=91;
				end
				if(in == 3) begin
					state<=1360;
					out<=92;
				end
				if(in == 4) begin
					state<=5249;
					out<=93;
				end
			end
			2118: begin
				if(in == 0) begin
					state<=2119;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=6008;
					out<=96;
				end
				if(in == 3) begin
					state<=121;
					out<=97;
				end
				if(in == 4) begin
					state<=4019;
					out<=98;
				end
			end
			2119: begin
				if(in == 0) begin
					state<=2120;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=6009;
					out<=101;
				end
				if(in == 3) begin
					state<=122;
					out<=102;
				end
				if(in == 4) begin
					state<=4020;
					out<=103;
				end
			end
			2120: begin
				if(in == 0) begin
					state<=2121;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=6010;
					out<=106;
				end
				if(in == 3) begin
					state<=123;
					out<=107;
				end
				if(in == 4) begin
					state<=4021;
					out<=108;
				end
			end
			2121: begin
				if(in == 0) begin
					state<=2122;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=6011;
					out<=111;
				end
				if(in == 3) begin
					state<=124;
					out<=112;
				end
				if(in == 4) begin
					state<=4022;
					out<=113;
				end
			end
			2122: begin
				if(in == 0) begin
					state<=2123;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=6012;
					out<=116;
				end
				if(in == 3) begin
					state<=125;
					out<=117;
				end
				if(in == 4) begin
					state<=4023;
					out<=118;
				end
			end
			2123: begin
				if(in == 0) begin
					state<=2124;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=6013;
					out<=121;
				end
				if(in == 3) begin
					state<=126;
					out<=122;
				end
				if(in == 4) begin
					state<=4024;
					out<=123;
				end
			end
			2124: begin
				if(in == 0) begin
					state<=2125;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=6014;
					out<=126;
				end
				if(in == 3) begin
					state<=127;
					out<=127;
				end
				if(in == 4) begin
					state<=4025;
					out<=128;
				end
			end
			2125: begin
				if(in == 0) begin
					state<=2126;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=6015;
					out<=131;
				end
				if(in == 3) begin
					state<=128;
					out<=132;
				end
				if(in == 4) begin
					state<=4026;
					out<=133;
				end
			end
			2126: begin
				if(in == 0) begin
					state<=2127;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=6016;
					out<=136;
				end
				if(in == 3) begin
					state<=129;
					out<=137;
				end
				if(in == 4) begin
					state<=4027;
					out<=138;
				end
			end
			2127: begin
				if(in == 0) begin
					state<=2128;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=6017;
					out<=141;
				end
				if(in == 3) begin
					state<=130;
					out<=142;
				end
				if(in == 4) begin
					state<=4028;
					out<=143;
				end
			end
			2128: begin
				if(in == 0) begin
					state<=2129;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=6018;
					out<=146;
				end
				if(in == 3) begin
					state<=131;
					out<=147;
				end
				if(in == 4) begin
					state<=4029;
					out<=148;
				end
			end
			2129: begin
				if(in == 0) begin
					state<=2130;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=6019;
					out<=151;
				end
				if(in == 3) begin
					state<=132;
					out<=152;
				end
				if(in == 4) begin
					state<=4030;
					out<=153;
				end
			end
			2130: begin
				if(in == 0) begin
					state<=2131;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=6020;
					out<=156;
				end
				if(in == 3) begin
					state<=133;
					out<=157;
				end
				if(in == 4) begin
					state<=4031;
					out<=158;
				end
			end
			2131: begin
				if(in == 0) begin
					state<=2132;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=6021;
					out<=161;
				end
				if(in == 3) begin
					state<=134;
					out<=162;
				end
				if(in == 4) begin
					state<=4032;
					out<=163;
				end
			end
			2132: begin
				if(in == 0) begin
					state<=2133;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=6022;
					out<=166;
				end
				if(in == 3) begin
					state<=135;
					out<=167;
				end
				if(in == 4) begin
					state<=4033;
					out<=168;
				end
			end
			2133: begin
				if(in == 0) begin
					state<=2134;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=6023;
					out<=171;
				end
				if(in == 3) begin
					state<=136;
					out<=172;
				end
				if(in == 4) begin
					state<=4034;
					out<=173;
				end
			end
			2134: begin
				if(in == 0) begin
					state<=2135;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=6024;
					out<=176;
				end
				if(in == 3) begin
					state<=137;
					out<=177;
				end
				if(in == 4) begin
					state<=4035;
					out<=178;
				end
			end
			2135: begin
				if(in == 0) begin
					state<=2136;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=6025;
					out<=181;
				end
				if(in == 3) begin
					state<=138;
					out<=182;
				end
				if(in == 4) begin
					state<=4036;
					out<=183;
				end
			end
			2136: begin
				if(in == 0) begin
					state<=2137;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=6026;
					out<=186;
				end
				if(in == 3) begin
					state<=139;
					out<=187;
				end
				if(in == 4) begin
					state<=4037;
					out<=188;
				end
			end
			2137: begin
				if(in == 0) begin
					state<=2138;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=6027;
					out<=191;
				end
				if(in == 3) begin
					state<=140;
					out<=192;
				end
				if(in == 4) begin
					state<=4038;
					out<=193;
				end
			end
			2138: begin
				if(in == 0) begin
					state<=2139;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=6028;
					out<=196;
				end
				if(in == 3) begin
					state<=141;
					out<=197;
				end
				if(in == 4) begin
					state<=4039;
					out<=198;
				end
			end
			2139: begin
				if(in == 0) begin
					state<=2140;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=6029;
					out<=201;
				end
				if(in == 3) begin
					state<=142;
					out<=202;
				end
				if(in == 4) begin
					state<=4040;
					out<=203;
				end
			end
			2140: begin
				if(in == 0) begin
					state<=2141;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=6030;
					out<=206;
				end
				if(in == 3) begin
					state<=143;
					out<=207;
				end
				if(in == 4) begin
					state<=4041;
					out<=208;
				end
			end
			2141: begin
				if(in == 0) begin
					state<=2142;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=6031;
					out<=211;
				end
				if(in == 3) begin
					state<=144;
					out<=212;
				end
				if(in == 4) begin
					state<=4042;
					out<=213;
				end
			end
			2142: begin
				if(in == 0) begin
					state<=2143;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=6032;
					out<=216;
				end
				if(in == 3) begin
					state<=145;
					out<=217;
				end
				if(in == 4) begin
					state<=4043;
					out<=218;
				end
			end
			2143: begin
				if(in == 0) begin
					state<=2144;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=6033;
					out<=221;
				end
				if(in == 3) begin
					state<=146;
					out<=222;
				end
				if(in == 4) begin
					state<=4044;
					out<=223;
				end
			end
			2144: begin
				if(in == 0) begin
					state<=2145;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=6034;
					out<=226;
				end
				if(in == 3) begin
					state<=147;
					out<=227;
				end
				if(in == 4) begin
					state<=4045;
					out<=228;
				end
			end
			2145: begin
				if(in == 0) begin
					state<=2146;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=6035;
					out<=231;
				end
				if(in == 3) begin
					state<=148;
					out<=232;
				end
				if(in == 4) begin
					state<=4046;
					out<=233;
				end
			end
			2146: begin
				if(in == 0) begin
					state<=2147;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=6036;
					out<=236;
				end
				if(in == 3) begin
					state<=149;
					out<=237;
				end
				if(in == 4) begin
					state<=4047;
					out<=238;
				end
			end
			2147: begin
				if(in == 0) begin
					state<=2148;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=6037;
					out<=241;
				end
				if(in == 3) begin
					state<=150;
					out<=242;
				end
				if(in == 4) begin
					state<=4048;
					out<=243;
				end
			end
			2148: begin
				if(in == 0) begin
					state<=2149;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=6038;
					out<=246;
				end
				if(in == 3) begin
					state<=151;
					out<=247;
				end
				if(in == 4) begin
					state<=4049;
					out<=248;
				end
			end
			2149: begin
				if(in == 0) begin
					state<=2150;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=6039;
					out<=251;
				end
				if(in == 3) begin
					state<=152;
					out<=252;
				end
				if(in == 4) begin
					state<=4050;
					out<=253;
				end
			end
			2150: begin
				if(in == 0) begin
					state<=2151;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=6040;
					out<=0;
				end
				if(in == 3) begin
					state<=153;
					out<=1;
				end
				if(in == 4) begin
					state<=4051;
					out<=2;
				end
			end
			2151: begin
				if(in == 0) begin
					state<=2152;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=6041;
					out<=5;
				end
				if(in == 3) begin
					state<=154;
					out<=6;
				end
				if(in == 4) begin
					state<=4052;
					out<=7;
				end
			end
			2152: begin
				if(in == 0) begin
					state<=2153;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=6042;
					out<=10;
				end
				if(in == 3) begin
					state<=155;
					out<=11;
				end
				if(in == 4) begin
					state<=4053;
					out<=12;
				end
			end
			2153: begin
				if(in == 0) begin
					state<=2154;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=6043;
					out<=15;
				end
				if(in == 3) begin
					state<=156;
					out<=16;
				end
				if(in == 4) begin
					state<=4054;
					out<=17;
				end
			end
			2154: begin
				if(in == 0) begin
					state<=2155;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=6044;
					out<=20;
				end
				if(in == 3) begin
					state<=157;
					out<=21;
				end
				if(in == 4) begin
					state<=4055;
					out<=22;
				end
			end
			2155: begin
				if(in == 0) begin
					state<=2156;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=6045;
					out<=25;
				end
				if(in == 3) begin
					state<=158;
					out<=26;
				end
				if(in == 4) begin
					state<=4056;
					out<=27;
				end
			end
			2156: begin
				if(in == 0) begin
					state<=2157;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=6046;
					out<=30;
				end
				if(in == 3) begin
					state<=159;
					out<=31;
				end
				if(in == 4) begin
					state<=4057;
					out<=32;
				end
			end
			2157: begin
				if(in == 0) begin
					state<=2158;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=6047;
					out<=35;
				end
				if(in == 3) begin
					state<=160;
					out<=36;
				end
				if(in == 4) begin
					state<=4058;
					out<=37;
				end
			end
			2158: begin
				if(in == 0) begin
					state<=2159;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=6048;
					out<=40;
				end
				if(in == 3) begin
					state<=161;
					out<=41;
				end
				if(in == 4) begin
					state<=4059;
					out<=42;
				end
			end
			2159: begin
				if(in == 0) begin
					state<=2160;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=6049;
					out<=45;
				end
				if(in == 3) begin
					state<=162;
					out<=46;
				end
				if(in == 4) begin
					state<=4060;
					out<=47;
				end
			end
			2160: begin
				if(in == 0) begin
					state<=2161;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=6050;
					out<=50;
				end
				if(in == 3) begin
					state<=163;
					out<=51;
				end
				if(in == 4) begin
					state<=4061;
					out<=52;
				end
			end
			2161: begin
				if(in == 0) begin
					state<=2162;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=6051;
					out<=55;
				end
				if(in == 3) begin
					state<=164;
					out<=56;
				end
				if(in == 4) begin
					state<=4062;
					out<=57;
				end
			end
			2162: begin
				if(in == 0) begin
					state<=2163;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=6052;
					out<=60;
				end
				if(in == 3) begin
					state<=165;
					out<=61;
				end
				if(in == 4) begin
					state<=4063;
					out<=62;
				end
			end
			2163: begin
				if(in == 0) begin
					state<=2164;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=6053;
					out<=65;
				end
				if(in == 3) begin
					state<=166;
					out<=66;
				end
				if(in == 4) begin
					state<=4064;
					out<=67;
				end
			end
			2164: begin
				if(in == 0) begin
					state<=2165;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=6054;
					out<=70;
				end
				if(in == 3) begin
					state<=167;
					out<=71;
				end
				if(in == 4) begin
					state<=4065;
					out<=72;
				end
			end
			2165: begin
				if(in == 0) begin
					state<=2166;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=6055;
					out<=75;
				end
				if(in == 3) begin
					state<=168;
					out<=76;
				end
				if(in == 4) begin
					state<=4066;
					out<=77;
				end
			end
			2166: begin
				if(in == 0) begin
					state<=2167;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=6056;
					out<=80;
				end
				if(in == 3) begin
					state<=169;
					out<=81;
				end
				if(in == 4) begin
					state<=4067;
					out<=82;
				end
			end
			2167: begin
				if(in == 0) begin
					state<=2168;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=6057;
					out<=85;
				end
				if(in == 3) begin
					state<=170;
					out<=86;
				end
				if(in == 4) begin
					state<=4068;
					out<=87;
				end
			end
			2168: begin
				if(in == 0) begin
					state<=2169;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=6058;
					out<=90;
				end
				if(in == 3) begin
					state<=171;
					out<=91;
				end
				if(in == 4) begin
					state<=4069;
					out<=92;
				end
			end
			2169: begin
				if(in == 0) begin
					state<=2170;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=6059;
					out<=95;
				end
				if(in == 3) begin
					state<=172;
					out<=96;
				end
				if(in == 4) begin
					state<=4070;
					out<=97;
				end
			end
			2170: begin
				if(in == 0) begin
					state<=2171;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=6060;
					out<=100;
				end
				if(in == 3) begin
					state<=173;
					out<=101;
				end
				if(in == 4) begin
					state<=4071;
					out<=102;
				end
			end
			2171: begin
				if(in == 0) begin
					state<=2172;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=6061;
					out<=105;
				end
				if(in == 3) begin
					state<=174;
					out<=106;
				end
				if(in == 4) begin
					state<=4072;
					out<=107;
				end
			end
			2172: begin
				if(in == 0) begin
					state<=2173;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=6062;
					out<=110;
				end
				if(in == 3) begin
					state<=175;
					out<=111;
				end
				if(in == 4) begin
					state<=4073;
					out<=112;
				end
			end
			2173: begin
				if(in == 0) begin
					state<=2174;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=6063;
					out<=115;
				end
				if(in == 3) begin
					state<=176;
					out<=116;
				end
				if(in == 4) begin
					state<=4074;
					out<=117;
				end
			end
			2174: begin
				if(in == 0) begin
					state<=2175;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=6064;
					out<=120;
				end
				if(in == 3) begin
					state<=177;
					out<=121;
				end
				if(in == 4) begin
					state<=4075;
					out<=122;
				end
			end
			2175: begin
				if(in == 0) begin
					state<=2176;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=6065;
					out<=125;
				end
				if(in == 3) begin
					state<=178;
					out<=126;
				end
				if(in == 4) begin
					state<=4076;
					out<=127;
				end
			end
			2176: begin
				if(in == 0) begin
					state<=2177;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=6066;
					out<=130;
				end
				if(in == 3) begin
					state<=179;
					out<=131;
				end
				if(in == 4) begin
					state<=4077;
					out<=132;
				end
			end
			2177: begin
				if(in == 0) begin
					state<=2178;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=6067;
					out<=135;
				end
				if(in == 3) begin
					state<=180;
					out<=136;
				end
				if(in == 4) begin
					state<=4078;
					out<=137;
				end
			end
			2178: begin
				if(in == 0) begin
					state<=2179;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=6068;
					out<=140;
				end
				if(in == 3) begin
					state<=181;
					out<=141;
				end
				if(in == 4) begin
					state<=4079;
					out<=142;
				end
			end
			2179: begin
				if(in == 0) begin
					state<=2180;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=6069;
					out<=145;
				end
				if(in == 3) begin
					state<=182;
					out<=146;
				end
				if(in == 4) begin
					state<=4080;
					out<=147;
				end
			end
			2180: begin
				if(in == 0) begin
					state<=2181;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=6070;
					out<=150;
				end
				if(in == 3) begin
					state<=183;
					out<=151;
				end
				if(in == 4) begin
					state<=4081;
					out<=152;
				end
			end
			2181: begin
				if(in == 0) begin
					state<=2182;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=6071;
					out<=155;
				end
				if(in == 3) begin
					state<=184;
					out<=156;
				end
				if(in == 4) begin
					state<=4082;
					out<=157;
				end
			end
			2182: begin
				if(in == 0) begin
					state<=2183;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=6072;
					out<=160;
				end
				if(in == 3) begin
					state<=185;
					out<=161;
				end
				if(in == 4) begin
					state<=4083;
					out<=162;
				end
			end
			2183: begin
				if(in == 0) begin
					state<=2184;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=6073;
					out<=165;
				end
				if(in == 3) begin
					state<=186;
					out<=166;
				end
				if(in == 4) begin
					state<=4084;
					out<=167;
				end
			end
			2184: begin
				if(in == 0) begin
					state<=2185;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=6074;
					out<=170;
				end
				if(in == 3) begin
					state<=187;
					out<=171;
				end
				if(in == 4) begin
					state<=4085;
					out<=172;
				end
			end
			2185: begin
				if(in == 0) begin
					state<=2186;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=6075;
					out<=175;
				end
				if(in == 3) begin
					state<=188;
					out<=176;
				end
				if(in == 4) begin
					state<=4086;
					out<=177;
				end
			end
			2186: begin
				if(in == 0) begin
					state<=3323;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=7212;
					out<=180;
				end
				if(in == 3) begin
					state<=1391;
					out<=181;
				end
				if(in == 4) begin
					state<=5280;
					out<=182;
				end
			end
			2187: begin
				if(in == 0) begin
					state<=2188;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=6077;
					out<=185;
				end
				if(in == 3) begin
					state<=190;
					out<=186;
				end
				if(in == 4) begin
					state<=4088;
					out<=187;
				end
			end
			2188: begin
				if(in == 0) begin
					state<=2189;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=6078;
					out<=190;
				end
				if(in == 3) begin
					state<=191;
					out<=191;
				end
				if(in == 4) begin
					state<=4089;
					out<=192;
				end
			end
			2189: begin
				if(in == 0) begin
					state<=2190;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=6079;
					out<=195;
				end
				if(in == 3) begin
					state<=192;
					out<=196;
				end
				if(in == 4) begin
					state<=4090;
					out<=197;
				end
			end
			2190: begin
				if(in == 0) begin
					state<=2191;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=6080;
					out<=200;
				end
				if(in == 3) begin
					state<=193;
					out<=201;
				end
				if(in == 4) begin
					state<=4091;
					out<=202;
				end
			end
			2191: begin
				if(in == 0) begin
					state<=2192;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=6081;
					out<=205;
				end
				if(in == 3) begin
					state<=194;
					out<=206;
				end
				if(in == 4) begin
					state<=4092;
					out<=207;
				end
			end
			2192: begin
				if(in == 0) begin
					state<=2193;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=6082;
					out<=210;
				end
				if(in == 3) begin
					state<=195;
					out<=211;
				end
				if(in == 4) begin
					state<=4093;
					out<=212;
				end
			end
			2193: begin
				if(in == 0) begin
					state<=2194;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=6083;
					out<=215;
				end
				if(in == 3) begin
					state<=196;
					out<=216;
				end
				if(in == 4) begin
					state<=4094;
					out<=217;
				end
			end
			2194: begin
				if(in == 0) begin
					state<=2195;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=6084;
					out<=220;
				end
				if(in == 3) begin
					state<=197;
					out<=221;
				end
				if(in == 4) begin
					state<=4095;
					out<=222;
				end
			end
			2195: begin
				if(in == 0) begin
					state<=2196;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=6085;
					out<=225;
				end
				if(in == 3) begin
					state<=198;
					out<=226;
				end
				if(in == 4) begin
					state<=4096;
					out<=227;
				end
			end
			2196: begin
				if(in == 0) begin
					state<=2197;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=6086;
					out<=230;
				end
				if(in == 3) begin
					state<=199;
					out<=231;
				end
				if(in == 4) begin
					state<=4097;
					out<=232;
				end
			end
			2197: begin
				if(in == 0) begin
					state<=2198;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=6087;
					out<=235;
				end
				if(in == 3) begin
					state<=200;
					out<=236;
				end
				if(in == 4) begin
					state<=4098;
					out<=237;
				end
			end
			2198: begin
				if(in == 0) begin
					state<=2199;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=6088;
					out<=240;
				end
				if(in == 3) begin
					state<=201;
					out<=241;
				end
				if(in == 4) begin
					state<=4099;
					out<=242;
				end
			end
			2199: begin
				if(in == 0) begin
					state<=2200;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=6089;
					out<=245;
				end
				if(in == 3) begin
					state<=202;
					out<=246;
				end
				if(in == 4) begin
					state<=4100;
					out<=247;
				end
			end
			2200: begin
				if(in == 0) begin
					state<=2201;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=6090;
					out<=250;
				end
				if(in == 3) begin
					state<=203;
					out<=251;
				end
				if(in == 4) begin
					state<=4101;
					out<=252;
				end
			end
			2201: begin
				if(in == 0) begin
					state<=2202;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=6091;
					out<=255;
				end
				if(in == 3) begin
					state<=204;
					out<=0;
				end
				if(in == 4) begin
					state<=4102;
					out<=1;
				end
			end
			2202: begin
				if(in == 0) begin
					state<=2203;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=6092;
					out<=4;
				end
				if(in == 3) begin
					state<=205;
					out<=5;
				end
				if(in == 4) begin
					state<=4103;
					out<=6;
				end
			end
			2203: begin
				if(in == 0) begin
					state<=2204;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=6093;
					out<=9;
				end
				if(in == 3) begin
					state<=206;
					out<=10;
				end
				if(in == 4) begin
					state<=4104;
					out<=11;
				end
			end
			2204: begin
				if(in == 0) begin
					state<=2205;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=6094;
					out<=14;
				end
				if(in == 3) begin
					state<=207;
					out<=15;
				end
				if(in == 4) begin
					state<=4105;
					out<=16;
				end
			end
			2205: begin
				if(in == 0) begin
					state<=2206;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=6095;
					out<=19;
				end
				if(in == 3) begin
					state<=208;
					out<=20;
				end
				if(in == 4) begin
					state<=4106;
					out<=21;
				end
			end
			2206: begin
				if(in == 0) begin
					state<=2207;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=6096;
					out<=24;
				end
				if(in == 3) begin
					state<=209;
					out<=25;
				end
				if(in == 4) begin
					state<=4107;
					out<=26;
				end
			end
			2207: begin
				if(in == 0) begin
					state<=2208;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=6097;
					out<=29;
				end
				if(in == 3) begin
					state<=210;
					out<=30;
				end
				if(in == 4) begin
					state<=4108;
					out<=31;
				end
			end
			2208: begin
				if(in == 0) begin
					state<=2209;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=6098;
					out<=34;
				end
				if(in == 3) begin
					state<=211;
					out<=35;
				end
				if(in == 4) begin
					state<=4109;
					out<=36;
				end
			end
			2209: begin
				if(in == 0) begin
					state<=2210;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=6099;
					out<=39;
				end
				if(in == 3) begin
					state<=212;
					out<=40;
				end
				if(in == 4) begin
					state<=4110;
					out<=41;
				end
			end
			2210: begin
				if(in == 0) begin
					state<=2211;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=6100;
					out<=44;
				end
				if(in == 3) begin
					state<=213;
					out<=45;
				end
				if(in == 4) begin
					state<=4111;
					out<=46;
				end
			end
			2211: begin
				if(in == 0) begin
					state<=2212;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=6101;
					out<=49;
				end
				if(in == 3) begin
					state<=214;
					out<=50;
				end
				if(in == 4) begin
					state<=4112;
					out<=51;
				end
			end
			2212: begin
				if(in == 0) begin
					state<=2213;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=6102;
					out<=54;
				end
				if(in == 3) begin
					state<=215;
					out<=55;
				end
				if(in == 4) begin
					state<=4113;
					out<=56;
				end
			end
			2213: begin
				if(in == 0) begin
					state<=2214;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=6103;
					out<=59;
				end
				if(in == 3) begin
					state<=216;
					out<=60;
				end
				if(in == 4) begin
					state<=4114;
					out<=61;
				end
			end
			2214: begin
				if(in == 0) begin
					state<=2215;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=6104;
					out<=64;
				end
				if(in == 3) begin
					state<=217;
					out<=65;
				end
				if(in == 4) begin
					state<=4115;
					out<=66;
				end
			end
			2215: begin
				if(in == 0) begin
					state<=2216;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=6105;
					out<=69;
				end
				if(in == 3) begin
					state<=218;
					out<=70;
				end
				if(in == 4) begin
					state<=4116;
					out<=71;
				end
			end
			2216: begin
				if(in == 0) begin
					state<=2217;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=6106;
					out<=74;
				end
				if(in == 3) begin
					state<=219;
					out<=75;
				end
				if(in == 4) begin
					state<=4117;
					out<=76;
				end
			end
			2217: begin
				if(in == 0) begin
					state<=2218;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=6107;
					out<=79;
				end
				if(in == 3) begin
					state<=220;
					out<=80;
				end
				if(in == 4) begin
					state<=4118;
					out<=81;
				end
			end
			2218: begin
				if(in == 0) begin
					state<=2219;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=6108;
					out<=84;
				end
				if(in == 3) begin
					state<=221;
					out<=85;
				end
				if(in == 4) begin
					state<=4119;
					out<=86;
				end
			end
			2219: begin
				if(in == 0) begin
					state<=2220;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=6109;
					out<=89;
				end
				if(in == 3) begin
					state<=222;
					out<=90;
				end
				if(in == 4) begin
					state<=4120;
					out<=91;
				end
			end
			2220: begin
				if(in == 0) begin
					state<=2221;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=6110;
					out<=94;
				end
				if(in == 3) begin
					state<=223;
					out<=95;
				end
				if(in == 4) begin
					state<=4121;
					out<=96;
				end
			end
			2221: begin
				if(in == 0) begin
					state<=2222;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=6111;
					out<=99;
				end
				if(in == 3) begin
					state<=224;
					out<=100;
				end
				if(in == 4) begin
					state<=4122;
					out<=101;
				end
			end
			2222: begin
				if(in == 0) begin
					state<=2223;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=6112;
					out<=104;
				end
				if(in == 3) begin
					state<=225;
					out<=105;
				end
				if(in == 4) begin
					state<=4123;
					out<=106;
				end
			end
			2223: begin
				if(in == 0) begin
					state<=2224;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=6113;
					out<=109;
				end
				if(in == 3) begin
					state<=226;
					out<=110;
				end
				if(in == 4) begin
					state<=4124;
					out<=111;
				end
			end
			2224: begin
				if(in == 0) begin
					state<=2225;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=6114;
					out<=114;
				end
				if(in == 3) begin
					state<=227;
					out<=115;
				end
				if(in == 4) begin
					state<=4125;
					out<=116;
				end
			end
			2225: begin
				if(in == 0) begin
					state<=2226;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=6115;
					out<=119;
				end
				if(in == 3) begin
					state<=228;
					out<=120;
				end
				if(in == 4) begin
					state<=4126;
					out<=121;
				end
			end
			2226: begin
				if(in == 0) begin
					state<=2227;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=6116;
					out<=124;
				end
				if(in == 3) begin
					state<=229;
					out<=125;
				end
				if(in == 4) begin
					state<=4127;
					out<=126;
				end
			end
			2227: begin
				if(in == 0) begin
					state<=2228;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=6117;
					out<=129;
				end
				if(in == 3) begin
					state<=230;
					out<=130;
				end
				if(in == 4) begin
					state<=4128;
					out<=131;
				end
			end
			2228: begin
				if(in == 0) begin
					state<=2229;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=6118;
					out<=134;
				end
				if(in == 3) begin
					state<=231;
					out<=135;
				end
				if(in == 4) begin
					state<=4129;
					out<=136;
				end
			end
			2229: begin
				if(in == 0) begin
					state<=2230;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=6119;
					out<=139;
				end
				if(in == 3) begin
					state<=232;
					out<=140;
				end
				if(in == 4) begin
					state<=4130;
					out<=141;
				end
			end
			2230: begin
				if(in == 0) begin
					state<=2231;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=6120;
					out<=144;
				end
				if(in == 3) begin
					state<=233;
					out<=145;
				end
				if(in == 4) begin
					state<=4131;
					out<=146;
				end
			end
			2231: begin
				if(in == 0) begin
					state<=2232;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=6121;
					out<=149;
				end
				if(in == 3) begin
					state<=234;
					out<=150;
				end
				if(in == 4) begin
					state<=4132;
					out<=151;
				end
			end
			2232: begin
				if(in == 0) begin
					state<=2233;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=6122;
					out<=154;
				end
				if(in == 3) begin
					state<=235;
					out<=155;
				end
				if(in == 4) begin
					state<=4133;
					out<=156;
				end
			end
			2233: begin
				if(in == 0) begin
					state<=2234;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=6123;
					out<=159;
				end
				if(in == 3) begin
					state<=236;
					out<=160;
				end
				if(in == 4) begin
					state<=4134;
					out<=161;
				end
			end
			2234: begin
				if(in == 0) begin
					state<=2235;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=6124;
					out<=164;
				end
				if(in == 3) begin
					state<=237;
					out<=165;
				end
				if(in == 4) begin
					state<=4135;
					out<=166;
				end
			end
			2235: begin
				if(in == 0) begin
					state<=2236;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=6125;
					out<=169;
				end
				if(in == 3) begin
					state<=238;
					out<=170;
				end
				if(in == 4) begin
					state<=4136;
					out<=171;
				end
			end
			2236: begin
				if(in == 0) begin
					state<=2237;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=6126;
					out<=174;
				end
				if(in == 3) begin
					state<=239;
					out<=175;
				end
				if(in == 4) begin
					state<=4137;
					out<=176;
				end
			end
			2237: begin
				if(in == 0) begin
					state<=2238;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=6127;
					out<=179;
				end
				if(in == 3) begin
					state<=240;
					out<=180;
				end
				if(in == 4) begin
					state<=4138;
					out<=181;
				end
			end
			2238: begin
				if(in == 0) begin
					state<=2239;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=6128;
					out<=184;
				end
				if(in == 3) begin
					state<=241;
					out<=185;
				end
				if(in == 4) begin
					state<=4139;
					out<=186;
				end
			end
			2239: begin
				if(in == 0) begin
					state<=2240;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=6129;
					out<=189;
				end
				if(in == 3) begin
					state<=242;
					out<=190;
				end
				if(in == 4) begin
					state<=4140;
					out<=191;
				end
			end
			2240: begin
				if(in == 0) begin
					state<=2241;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=6130;
					out<=194;
				end
				if(in == 3) begin
					state<=243;
					out<=195;
				end
				if(in == 4) begin
					state<=4141;
					out<=196;
				end
			end
			2241: begin
				if(in == 0) begin
					state<=2242;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=6131;
					out<=199;
				end
				if(in == 3) begin
					state<=244;
					out<=200;
				end
				if(in == 4) begin
					state<=4142;
					out<=201;
				end
			end
			2242: begin
				if(in == 0) begin
					state<=2243;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=6132;
					out<=204;
				end
				if(in == 3) begin
					state<=245;
					out<=205;
				end
				if(in == 4) begin
					state<=4143;
					out<=206;
				end
			end
			2243: begin
				if(in == 0) begin
					state<=2244;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=6133;
					out<=209;
				end
				if(in == 3) begin
					state<=246;
					out<=210;
				end
				if(in == 4) begin
					state<=4144;
					out<=211;
				end
			end
			2244: begin
				if(in == 0) begin
					state<=2245;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=6134;
					out<=214;
				end
				if(in == 3) begin
					state<=247;
					out<=215;
				end
				if(in == 4) begin
					state<=4145;
					out<=216;
				end
			end
			2245: begin
				if(in == 0) begin
					state<=2246;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=6135;
					out<=219;
				end
				if(in == 3) begin
					state<=248;
					out<=220;
				end
				if(in == 4) begin
					state<=4146;
					out<=221;
				end
			end
			2246: begin
				if(in == 0) begin
					state<=2247;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=6136;
					out<=224;
				end
				if(in == 3) begin
					state<=249;
					out<=225;
				end
				if(in == 4) begin
					state<=4147;
					out<=226;
				end
			end
			2247: begin
				if(in == 0) begin
					state<=2248;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=6137;
					out<=229;
				end
				if(in == 3) begin
					state<=250;
					out<=230;
				end
				if(in == 4) begin
					state<=4148;
					out<=231;
				end
			end
			2248: begin
				if(in == 0) begin
					state<=2249;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=6138;
					out<=234;
				end
				if(in == 3) begin
					state<=251;
					out<=235;
				end
				if(in == 4) begin
					state<=4149;
					out<=236;
				end
			end
			2249: begin
				if(in == 0) begin
					state<=2250;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=6139;
					out<=239;
				end
				if(in == 3) begin
					state<=252;
					out<=240;
				end
				if(in == 4) begin
					state<=4150;
					out<=241;
				end
			end
			2250: begin
				if(in == 0) begin
					state<=2251;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=6140;
					out<=244;
				end
				if(in == 3) begin
					state<=253;
					out<=245;
				end
				if(in == 4) begin
					state<=4151;
					out<=246;
				end
			end
			2251: begin
				if(in == 0) begin
					state<=2252;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=6141;
					out<=249;
				end
				if(in == 3) begin
					state<=254;
					out<=250;
				end
				if(in == 4) begin
					state<=4152;
					out<=251;
				end
			end
			2252: begin
				if(in == 0) begin
					state<=2253;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=6142;
					out<=254;
				end
				if(in == 3) begin
					state<=255;
					out<=255;
				end
				if(in == 4) begin
					state<=4153;
					out<=0;
				end
			end
			2253: begin
				if(in == 0) begin
					state<=2254;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=6143;
					out<=3;
				end
				if(in == 3) begin
					state<=256;
					out<=4;
				end
				if(in == 4) begin
					state<=4154;
					out<=5;
				end
			end
			2254: begin
				if(in == 0) begin
					state<=2255;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=6144;
					out<=8;
				end
				if(in == 3) begin
					state<=257;
					out<=9;
				end
				if(in == 4) begin
					state<=4155;
					out<=10;
				end
			end
			2255: begin
				if(in == 0) begin
					state<=3354;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=7243;
					out<=13;
				end
				if(in == 3) begin
					state<=1422;
					out<=14;
				end
				if(in == 4) begin
					state<=5311;
					out<=15;
				end
			end
			2256: begin
				if(in == 0) begin
					state<=2257;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=6146;
					out<=18;
				end
				if(in == 3) begin
					state<=259;
					out<=19;
				end
				if(in == 4) begin
					state<=4157;
					out<=20;
				end
			end
			2257: begin
				if(in == 0) begin
					state<=2258;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=6147;
					out<=23;
				end
				if(in == 3) begin
					state<=260;
					out<=24;
				end
				if(in == 4) begin
					state<=4158;
					out<=25;
				end
			end
			2258: begin
				if(in == 0) begin
					state<=2259;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=6148;
					out<=28;
				end
				if(in == 3) begin
					state<=261;
					out<=29;
				end
				if(in == 4) begin
					state<=4159;
					out<=30;
				end
			end
			2259: begin
				if(in == 0) begin
					state<=2260;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=6149;
					out<=33;
				end
				if(in == 3) begin
					state<=262;
					out<=34;
				end
				if(in == 4) begin
					state<=4160;
					out<=35;
				end
			end
			2260: begin
				if(in == 0) begin
					state<=2261;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=6150;
					out<=38;
				end
				if(in == 3) begin
					state<=263;
					out<=39;
				end
				if(in == 4) begin
					state<=4161;
					out<=40;
				end
			end
			2261: begin
				if(in == 0) begin
					state<=2262;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=6151;
					out<=43;
				end
				if(in == 3) begin
					state<=264;
					out<=44;
				end
				if(in == 4) begin
					state<=4162;
					out<=45;
				end
			end
			2262: begin
				if(in == 0) begin
					state<=2263;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=6152;
					out<=48;
				end
				if(in == 3) begin
					state<=265;
					out<=49;
				end
				if(in == 4) begin
					state<=4163;
					out<=50;
				end
			end
			2263: begin
				if(in == 0) begin
					state<=2264;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=6153;
					out<=53;
				end
				if(in == 3) begin
					state<=266;
					out<=54;
				end
				if(in == 4) begin
					state<=4164;
					out<=55;
				end
			end
			2264: begin
				if(in == 0) begin
					state<=2265;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=6154;
					out<=58;
				end
				if(in == 3) begin
					state<=267;
					out<=59;
				end
				if(in == 4) begin
					state<=4165;
					out<=60;
				end
			end
			2265: begin
				if(in == 0) begin
					state<=2266;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=6155;
					out<=63;
				end
				if(in == 3) begin
					state<=268;
					out<=64;
				end
				if(in == 4) begin
					state<=4166;
					out<=65;
				end
			end
			2266: begin
				if(in == 0) begin
					state<=2267;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=6156;
					out<=68;
				end
				if(in == 3) begin
					state<=269;
					out<=69;
				end
				if(in == 4) begin
					state<=4167;
					out<=70;
				end
			end
			2267: begin
				if(in == 0) begin
					state<=2268;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=6157;
					out<=73;
				end
				if(in == 3) begin
					state<=270;
					out<=74;
				end
				if(in == 4) begin
					state<=4168;
					out<=75;
				end
			end
			2268: begin
				if(in == 0) begin
					state<=2269;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=6158;
					out<=78;
				end
				if(in == 3) begin
					state<=271;
					out<=79;
				end
				if(in == 4) begin
					state<=4169;
					out<=80;
				end
			end
			2269: begin
				if(in == 0) begin
					state<=2270;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=6159;
					out<=83;
				end
				if(in == 3) begin
					state<=272;
					out<=84;
				end
				if(in == 4) begin
					state<=4170;
					out<=85;
				end
			end
			2270: begin
				if(in == 0) begin
					state<=2271;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=6160;
					out<=88;
				end
				if(in == 3) begin
					state<=273;
					out<=89;
				end
				if(in == 4) begin
					state<=4171;
					out<=90;
				end
			end
			2271: begin
				if(in == 0) begin
					state<=2272;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=6161;
					out<=93;
				end
				if(in == 3) begin
					state<=274;
					out<=94;
				end
				if(in == 4) begin
					state<=4172;
					out<=95;
				end
			end
			2272: begin
				if(in == 0) begin
					state<=2273;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=6162;
					out<=98;
				end
				if(in == 3) begin
					state<=275;
					out<=99;
				end
				if(in == 4) begin
					state<=4173;
					out<=100;
				end
			end
			2273: begin
				if(in == 0) begin
					state<=2274;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=6163;
					out<=103;
				end
				if(in == 3) begin
					state<=276;
					out<=104;
				end
				if(in == 4) begin
					state<=4174;
					out<=105;
				end
			end
			2274: begin
				if(in == 0) begin
					state<=2275;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=6164;
					out<=108;
				end
				if(in == 3) begin
					state<=277;
					out<=109;
				end
				if(in == 4) begin
					state<=4175;
					out<=110;
				end
			end
			2275: begin
				if(in == 0) begin
					state<=2276;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=6165;
					out<=113;
				end
				if(in == 3) begin
					state<=278;
					out<=114;
				end
				if(in == 4) begin
					state<=4176;
					out<=115;
				end
			end
			2276: begin
				if(in == 0) begin
					state<=2277;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=6166;
					out<=118;
				end
				if(in == 3) begin
					state<=279;
					out<=119;
				end
				if(in == 4) begin
					state<=4177;
					out<=120;
				end
			end
			2277: begin
				if(in == 0) begin
					state<=2278;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=6167;
					out<=123;
				end
				if(in == 3) begin
					state<=280;
					out<=124;
				end
				if(in == 4) begin
					state<=4178;
					out<=125;
				end
			end
			2278: begin
				if(in == 0) begin
					state<=2279;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=6168;
					out<=128;
				end
				if(in == 3) begin
					state<=281;
					out<=129;
				end
				if(in == 4) begin
					state<=4179;
					out<=130;
				end
			end
			2279: begin
				if(in == 0) begin
					state<=2280;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=6169;
					out<=133;
				end
				if(in == 3) begin
					state<=282;
					out<=134;
				end
				if(in == 4) begin
					state<=4180;
					out<=135;
				end
			end
			2280: begin
				if(in == 0) begin
					state<=2281;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=6170;
					out<=138;
				end
				if(in == 3) begin
					state<=283;
					out<=139;
				end
				if(in == 4) begin
					state<=4181;
					out<=140;
				end
			end
			2281: begin
				if(in == 0) begin
					state<=2282;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=6171;
					out<=143;
				end
				if(in == 3) begin
					state<=284;
					out<=144;
				end
				if(in == 4) begin
					state<=4182;
					out<=145;
				end
			end
			2282: begin
				if(in == 0) begin
					state<=2283;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=6172;
					out<=148;
				end
				if(in == 3) begin
					state<=285;
					out<=149;
				end
				if(in == 4) begin
					state<=4183;
					out<=150;
				end
			end
			2283: begin
				if(in == 0) begin
					state<=2284;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=6173;
					out<=153;
				end
				if(in == 3) begin
					state<=286;
					out<=154;
				end
				if(in == 4) begin
					state<=4184;
					out<=155;
				end
			end
			2284: begin
				if(in == 0) begin
					state<=2285;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=6174;
					out<=158;
				end
				if(in == 3) begin
					state<=287;
					out<=159;
				end
				if(in == 4) begin
					state<=4185;
					out<=160;
				end
			end
			2285: begin
				if(in == 0) begin
					state<=2286;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=6175;
					out<=163;
				end
				if(in == 3) begin
					state<=288;
					out<=164;
				end
				if(in == 4) begin
					state<=4186;
					out<=165;
				end
			end
			2286: begin
				if(in == 0) begin
					state<=2287;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=6176;
					out<=168;
				end
				if(in == 3) begin
					state<=289;
					out<=169;
				end
				if(in == 4) begin
					state<=4187;
					out<=170;
				end
			end
			2287: begin
				if(in == 0) begin
					state<=2288;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=6177;
					out<=173;
				end
				if(in == 3) begin
					state<=290;
					out<=174;
				end
				if(in == 4) begin
					state<=4188;
					out<=175;
				end
			end
			2288: begin
				if(in == 0) begin
					state<=2289;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=6178;
					out<=178;
				end
				if(in == 3) begin
					state<=291;
					out<=179;
				end
				if(in == 4) begin
					state<=4189;
					out<=180;
				end
			end
			2289: begin
				if(in == 0) begin
					state<=2290;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=6179;
					out<=183;
				end
				if(in == 3) begin
					state<=292;
					out<=184;
				end
				if(in == 4) begin
					state<=4190;
					out<=185;
				end
			end
			2290: begin
				if(in == 0) begin
					state<=2291;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=6180;
					out<=188;
				end
				if(in == 3) begin
					state<=293;
					out<=189;
				end
				if(in == 4) begin
					state<=4191;
					out<=190;
				end
			end
			2291: begin
				if(in == 0) begin
					state<=2292;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=6181;
					out<=193;
				end
				if(in == 3) begin
					state<=294;
					out<=194;
				end
				if(in == 4) begin
					state<=4192;
					out<=195;
				end
			end
			2292: begin
				if(in == 0) begin
					state<=2293;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=6182;
					out<=198;
				end
				if(in == 3) begin
					state<=295;
					out<=199;
				end
				if(in == 4) begin
					state<=4193;
					out<=200;
				end
			end
			2293: begin
				if(in == 0) begin
					state<=2294;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=6183;
					out<=203;
				end
				if(in == 3) begin
					state<=296;
					out<=204;
				end
				if(in == 4) begin
					state<=4194;
					out<=205;
				end
			end
			2294: begin
				if(in == 0) begin
					state<=2295;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=6184;
					out<=208;
				end
				if(in == 3) begin
					state<=297;
					out<=209;
				end
				if(in == 4) begin
					state<=4195;
					out<=210;
				end
			end
			2295: begin
				if(in == 0) begin
					state<=2296;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=6185;
					out<=213;
				end
				if(in == 3) begin
					state<=298;
					out<=214;
				end
				if(in == 4) begin
					state<=4196;
					out<=215;
				end
			end
			2296: begin
				if(in == 0) begin
					state<=2297;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=6186;
					out<=218;
				end
				if(in == 3) begin
					state<=299;
					out<=219;
				end
				if(in == 4) begin
					state<=4197;
					out<=220;
				end
			end
			2297: begin
				if(in == 0) begin
					state<=2298;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=6187;
					out<=223;
				end
				if(in == 3) begin
					state<=300;
					out<=224;
				end
				if(in == 4) begin
					state<=4198;
					out<=225;
				end
			end
			2298: begin
				if(in == 0) begin
					state<=2299;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=6188;
					out<=228;
				end
				if(in == 3) begin
					state<=301;
					out<=229;
				end
				if(in == 4) begin
					state<=4199;
					out<=230;
				end
			end
			2299: begin
				if(in == 0) begin
					state<=2300;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=6189;
					out<=233;
				end
				if(in == 3) begin
					state<=302;
					out<=234;
				end
				if(in == 4) begin
					state<=4200;
					out<=235;
				end
			end
			2300: begin
				if(in == 0) begin
					state<=2301;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=6190;
					out<=238;
				end
				if(in == 3) begin
					state<=303;
					out<=239;
				end
				if(in == 4) begin
					state<=4201;
					out<=240;
				end
			end
			2301: begin
				if(in == 0) begin
					state<=2302;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=6191;
					out<=243;
				end
				if(in == 3) begin
					state<=304;
					out<=244;
				end
				if(in == 4) begin
					state<=4202;
					out<=245;
				end
			end
			2302: begin
				if(in == 0) begin
					state<=2303;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=6192;
					out<=248;
				end
				if(in == 3) begin
					state<=305;
					out<=249;
				end
				if(in == 4) begin
					state<=4203;
					out<=250;
				end
			end
			2303: begin
				if(in == 0) begin
					state<=2304;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=6193;
					out<=253;
				end
				if(in == 3) begin
					state<=306;
					out<=254;
				end
				if(in == 4) begin
					state<=4204;
					out<=255;
				end
			end
			2304: begin
				if(in == 0) begin
					state<=2305;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=6194;
					out<=2;
				end
				if(in == 3) begin
					state<=307;
					out<=3;
				end
				if(in == 4) begin
					state<=4205;
					out<=4;
				end
			end
			2305: begin
				if(in == 0) begin
					state<=2306;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=6195;
					out<=7;
				end
				if(in == 3) begin
					state<=308;
					out<=8;
				end
				if(in == 4) begin
					state<=4206;
					out<=9;
				end
			end
			2306: begin
				if(in == 0) begin
					state<=2307;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=6196;
					out<=12;
				end
				if(in == 3) begin
					state<=309;
					out<=13;
				end
				if(in == 4) begin
					state<=4207;
					out<=14;
				end
			end
			2307: begin
				if(in == 0) begin
					state<=2308;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=6197;
					out<=17;
				end
				if(in == 3) begin
					state<=310;
					out<=18;
				end
				if(in == 4) begin
					state<=4208;
					out<=19;
				end
			end
			2308: begin
				if(in == 0) begin
					state<=2309;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=6198;
					out<=22;
				end
				if(in == 3) begin
					state<=311;
					out<=23;
				end
				if(in == 4) begin
					state<=4209;
					out<=24;
				end
			end
			2309: begin
				if(in == 0) begin
					state<=2310;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=6199;
					out<=27;
				end
				if(in == 3) begin
					state<=312;
					out<=28;
				end
				if(in == 4) begin
					state<=4210;
					out<=29;
				end
			end
			2310: begin
				if(in == 0) begin
					state<=2311;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=6200;
					out<=32;
				end
				if(in == 3) begin
					state<=313;
					out<=33;
				end
				if(in == 4) begin
					state<=4211;
					out<=34;
				end
			end
			2311: begin
				if(in == 0) begin
					state<=2312;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=6201;
					out<=37;
				end
				if(in == 3) begin
					state<=314;
					out<=38;
				end
				if(in == 4) begin
					state<=4212;
					out<=39;
				end
			end
			2312: begin
				if(in == 0) begin
					state<=2313;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=6202;
					out<=42;
				end
				if(in == 3) begin
					state<=315;
					out<=43;
				end
				if(in == 4) begin
					state<=4213;
					out<=44;
				end
			end
			2313: begin
				if(in == 0) begin
					state<=2314;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=6203;
					out<=47;
				end
				if(in == 3) begin
					state<=316;
					out<=48;
				end
				if(in == 4) begin
					state<=4214;
					out<=49;
				end
			end
			2314: begin
				if(in == 0) begin
					state<=2315;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=6204;
					out<=52;
				end
				if(in == 3) begin
					state<=317;
					out<=53;
				end
				if(in == 4) begin
					state<=4215;
					out<=54;
				end
			end
			2315: begin
				if(in == 0) begin
					state<=2316;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=6205;
					out<=57;
				end
				if(in == 3) begin
					state<=318;
					out<=58;
				end
				if(in == 4) begin
					state<=4216;
					out<=59;
				end
			end
			2316: begin
				if(in == 0) begin
					state<=2317;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=6206;
					out<=62;
				end
				if(in == 3) begin
					state<=319;
					out<=63;
				end
				if(in == 4) begin
					state<=4217;
					out<=64;
				end
			end
			2317: begin
				if(in == 0) begin
					state<=2318;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=6207;
					out<=67;
				end
				if(in == 3) begin
					state<=320;
					out<=68;
				end
				if(in == 4) begin
					state<=4218;
					out<=69;
				end
			end
			2318: begin
				if(in == 0) begin
					state<=2319;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=6208;
					out<=72;
				end
				if(in == 3) begin
					state<=321;
					out<=73;
				end
				if(in == 4) begin
					state<=4219;
					out<=74;
				end
			end
			2319: begin
				if(in == 0) begin
					state<=2320;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=6209;
					out<=77;
				end
				if(in == 3) begin
					state<=322;
					out<=78;
				end
				if(in == 4) begin
					state<=4220;
					out<=79;
				end
			end
			2320: begin
				if(in == 0) begin
					state<=2321;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=6210;
					out<=82;
				end
				if(in == 3) begin
					state<=323;
					out<=83;
				end
				if(in == 4) begin
					state<=4221;
					out<=84;
				end
			end
			2321: begin
				if(in == 0) begin
					state<=2322;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=6211;
					out<=87;
				end
				if(in == 3) begin
					state<=324;
					out<=88;
				end
				if(in == 4) begin
					state<=4222;
					out<=89;
				end
			end
			2322: begin
				if(in == 0) begin
					state<=2323;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=6212;
					out<=92;
				end
				if(in == 3) begin
					state<=325;
					out<=93;
				end
				if(in == 4) begin
					state<=4223;
					out<=94;
				end
			end
			2323: begin
				if(in == 0) begin
					state<=2324;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=6213;
					out<=97;
				end
				if(in == 3) begin
					state<=326;
					out<=98;
				end
				if(in == 4) begin
					state<=4224;
					out<=99;
				end
			end
			2324: begin
				if(in == 0) begin
					state<=2898;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=6787;
					out<=102;
				end
				if(in == 3) begin
					state<=1453;
					out<=103;
				end
				if(in == 4) begin
					state<=5342;
					out<=104;
				end
			end
			2325: begin
				if(in == 0) begin
					state<=2326;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=6215;
					out<=107;
				end
				if(in == 3) begin
					state<=328;
					out<=108;
				end
				if(in == 4) begin
					state<=4226;
					out<=109;
				end
			end
			2326: begin
				if(in == 0) begin
					state<=2327;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=6216;
					out<=112;
				end
				if(in == 3) begin
					state<=329;
					out<=113;
				end
				if(in == 4) begin
					state<=4227;
					out<=114;
				end
			end
			2327: begin
				if(in == 0) begin
					state<=2328;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=6217;
					out<=117;
				end
				if(in == 3) begin
					state<=330;
					out<=118;
				end
				if(in == 4) begin
					state<=4228;
					out<=119;
				end
			end
			2328: begin
				if(in == 0) begin
					state<=2329;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=6218;
					out<=122;
				end
				if(in == 3) begin
					state<=331;
					out<=123;
				end
				if(in == 4) begin
					state<=4229;
					out<=124;
				end
			end
			2329: begin
				if(in == 0) begin
					state<=2330;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=6219;
					out<=127;
				end
				if(in == 3) begin
					state<=332;
					out<=128;
				end
				if(in == 4) begin
					state<=4230;
					out<=129;
				end
			end
			2330: begin
				if(in == 0) begin
					state<=2331;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=6220;
					out<=132;
				end
				if(in == 3) begin
					state<=333;
					out<=133;
				end
				if(in == 4) begin
					state<=4231;
					out<=134;
				end
			end
			2331: begin
				if(in == 0) begin
					state<=2332;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=6221;
					out<=137;
				end
				if(in == 3) begin
					state<=334;
					out<=138;
				end
				if(in == 4) begin
					state<=4232;
					out<=139;
				end
			end
			2332: begin
				if(in == 0) begin
					state<=2333;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=6222;
					out<=142;
				end
				if(in == 3) begin
					state<=335;
					out<=143;
				end
				if(in == 4) begin
					state<=4233;
					out<=144;
				end
			end
			2333: begin
				if(in == 0) begin
					state<=2334;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=6223;
					out<=147;
				end
				if(in == 3) begin
					state<=336;
					out<=148;
				end
				if(in == 4) begin
					state<=4234;
					out<=149;
				end
			end
			2334: begin
				if(in == 0) begin
					state<=2335;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=6224;
					out<=152;
				end
				if(in == 3) begin
					state<=337;
					out<=153;
				end
				if(in == 4) begin
					state<=4235;
					out<=154;
				end
			end
			2335: begin
				if(in == 0) begin
					state<=2336;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=6225;
					out<=157;
				end
				if(in == 3) begin
					state<=338;
					out<=158;
				end
				if(in == 4) begin
					state<=4236;
					out<=159;
				end
			end
			2336: begin
				if(in == 0) begin
					state<=2337;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=6226;
					out<=162;
				end
				if(in == 3) begin
					state<=339;
					out<=163;
				end
				if(in == 4) begin
					state<=4237;
					out<=164;
				end
			end
			2337: begin
				if(in == 0) begin
					state<=2338;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=6227;
					out<=167;
				end
				if(in == 3) begin
					state<=340;
					out<=168;
				end
				if(in == 4) begin
					state<=4238;
					out<=169;
				end
			end
			2338: begin
				if(in == 0) begin
					state<=2339;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=6228;
					out<=172;
				end
				if(in == 3) begin
					state<=341;
					out<=173;
				end
				if(in == 4) begin
					state<=4239;
					out<=174;
				end
			end
			2339: begin
				if(in == 0) begin
					state<=2340;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=6229;
					out<=177;
				end
				if(in == 3) begin
					state<=342;
					out<=178;
				end
				if(in == 4) begin
					state<=4240;
					out<=179;
				end
			end
			2340: begin
				if(in == 0) begin
					state<=2341;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=6230;
					out<=182;
				end
				if(in == 3) begin
					state<=343;
					out<=183;
				end
				if(in == 4) begin
					state<=4241;
					out<=184;
				end
			end
			2341: begin
				if(in == 0) begin
					state<=2342;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=6231;
					out<=187;
				end
				if(in == 3) begin
					state<=344;
					out<=188;
				end
				if(in == 4) begin
					state<=4242;
					out<=189;
				end
			end
			2342: begin
				if(in == 0) begin
					state<=2343;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=6232;
					out<=192;
				end
				if(in == 3) begin
					state<=345;
					out<=193;
				end
				if(in == 4) begin
					state<=4243;
					out<=194;
				end
			end
			2343: begin
				if(in == 0) begin
					state<=2344;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=6233;
					out<=197;
				end
				if(in == 3) begin
					state<=346;
					out<=198;
				end
				if(in == 4) begin
					state<=4244;
					out<=199;
				end
			end
			2344: begin
				if(in == 0) begin
					state<=2345;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=6234;
					out<=202;
				end
				if(in == 3) begin
					state<=347;
					out<=203;
				end
				if(in == 4) begin
					state<=4245;
					out<=204;
				end
			end
			2345: begin
				if(in == 0) begin
					state<=2346;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=6235;
					out<=207;
				end
				if(in == 3) begin
					state<=348;
					out<=208;
				end
				if(in == 4) begin
					state<=4246;
					out<=209;
				end
			end
			2346: begin
				if(in == 0) begin
					state<=2347;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=6236;
					out<=212;
				end
				if(in == 3) begin
					state<=349;
					out<=213;
				end
				if(in == 4) begin
					state<=4247;
					out<=214;
				end
			end
			2347: begin
				if(in == 0) begin
					state<=2348;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=6237;
					out<=217;
				end
				if(in == 3) begin
					state<=350;
					out<=218;
				end
				if(in == 4) begin
					state<=4248;
					out<=219;
				end
			end
			2348: begin
				if(in == 0) begin
					state<=2349;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=6238;
					out<=222;
				end
				if(in == 3) begin
					state<=351;
					out<=223;
				end
				if(in == 4) begin
					state<=4249;
					out<=224;
				end
			end
			2349: begin
				if(in == 0) begin
					state<=2350;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=6239;
					out<=227;
				end
				if(in == 3) begin
					state<=352;
					out<=228;
				end
				if(in == 4) begin
					state<=4250;
					out<=229;
				end
			end
			2350: begin
				if(in == 0) begin
					state<=2351;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=6240;
					out<=232;
				end
				if(in == 3) begin
					state<=353;
					out<=233;
				end
				if(in == 4) begin
					state<=4251;
					out<=234;
				end
			end
			2351: begin
				if(in == 0) begin
					state<=2352;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=6241;
					out<=237;
				end
				if(in == 3) begin
					state<=354;
					out<=238;
				end
				if(in == 4) begin
					state<=4252;
					out<=239;
				end
			end
			2352: begin
				if(in == 0) begin
					state<=2353;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=6242;
					out<=242;
				end
				if(in == 3) begin
					state<=355;
					out<=243;
				end
				if(in == 4) begin
					state<=4253;
					out<=244;
				end
			end
			2353: begin
				if(in == 0) begin
					state<=2354;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=6243;
					out<=247;
				end
				if(in == 3) begin
					state<=356;
					out<=248;
				end
				if(in == 4) begin
					state<=4254;
					out<=249;
				end
			end
			2354: begin
				if(in == 0) begin
					state<=2355;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=6244;
					out<=252;
				end
				if(in == 3) begin
					state<=357;
					out<=253;
				end
				if(in == 4) begin
					state<=4255;
					out<=254;
				end
			end
			2355: begin
				if(in == 0) begin
					state<=2356;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=6245;
					out<=1;
				end
				if(in == 3) begin
					state<=358;
					out<=2;
				end
				if(in == 4) begin
					state<=4256;
					out<=3;
				end
			end
			2356: begin
				if(in == 0) begin
					state<=2357;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=6246;
					out<=6;
				end
				if(in == 3) begin
					state<=359;
					out<=7;
				end
				if(in == 4) begin
					state<=4257;
					out<=8;
				end
			end
			2357: begin
				if(in == 0) begin
					state<=2358;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=6247;
					out<=11;
				end
				if(in == 3) begin
					state<=360;
					out<=12;
				end
				if(in == 4) begin
					state<=4258;
					out<=13;
				end
			end
			2358: begin
				if(in == 0) begin
					state<=2359;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=6248;
					out<=16;
				end
				if(in == 3) begin
					state<=361;
					out<=17;
				end
				if(in == 4) begin
					state<=4259;
					out<=18;
				end
			end
			2359: begin
				if(in == 0) begin
					state<=2360;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=6249;
					out<=21;
				end
				if(in == 3) begin
					state<=362;
					out<=22;
				end
				if(in == 4) begin
					state<=4260;
					out<=23;
				end
			end
			2360: begin
				if(in == 0) begin
					state<=2361;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=6250;
					out<=26;
				end
				if(in == 3) begin
					state<=363;
					out<=27;
				end
				if(in == 4) begin
					state<=4261;
					out<=28;
				end
			end
			2361: begin
				if(in == 0) begin
					state<=2362;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=6251;
					out<=31;
				end
				if(in == 3) begin
					state<=364;
					out<=32;
				end
				if(in == 4) begin
					state<=4262;
					out<=33;
				end
			end
			2362: begin
				if(in == 0) begin
					state<=2363;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=6252;
					out<=36;
				end
				if(in == 3) begin
					state<=365;
					out<=37;
				end
				if(in == 4) begin
					state<=4263;
					out<=38;
				end
			end
			2363: begin
				if(in == 0) begin
					state<=2364;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=6253;
					out<=41;
				end
				if(in == 3) begin
					state<=366;
					out<=42;
				end
				if(in == 4) begin
					state<=4264;
					out<=43;
				end
			end
			2364: begin
				if(in == 0) begin
					state<=2365;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=6254;
					out<=46;
				end
				if(in == 3) begin
					state<=367;
					out<=47;
				end
				if(in == 4) begin
					state<=4265;
					out<=48;
				end
			end
			2365: begin
				if(in == 0) begin
					state<=2366;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=6255;
					out<=51;
				end
				if(in == 3) begin
					state<=368;
					out<=52;
				end
				if(in == 4) begin
					state<=4266;
					out<=53;
				end
			end
			2366: begin
				if(in == 0) begin
					state<=2367;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=6256;
					out<=56;
				end
				if(in == 3) begin
					state<=369;
					out<=57;
				end
				if(in == 4) begin
					state<=4267;
					out<=58;
				end
			end
			2367: begin
				if(in == 0) begin
					state<=2368;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=6257;
					out<=61;
				end
				if(in == 3) begin
					state<=370;
					out<=62;
				end
				if(in == 4) begin
					state<=4268;
					out<=63;
				end
			end
			2368: begin
				if(in == 0) begin
					state<=2369;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=6258;
					out<=66;
				end
				if(in == 3) begin
					state<=371;
					out<=67;
				end
				if(in == 4) begin
					state<=4269;
					out<=68;
				end
			end
			2369: begin
				if(in == 0) begin
					state<=2370;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=6259;
					out<=71;
				end
				if(in == 3) begin
					state<=372;
					out<=72;
				end
				if(in == 4) begin
					state<=4270;
					out<=73;
				end
			end
			2370: begin
				if(in == 0) begin
					state<=2371;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=6260;
					out<=76;
				end
				if(in == 3) begin
					state<=373;
					out<=77;
				end
				if(in == 4) begin
					state<=4271;
					out<=78;
				end
			end
			2371: begin
				if(in == 0) begin
					state<=2372;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=6261;
					out<=81;
				end
				if(in == 3) begin
					state<=374;
					out<=82;
				end
				if(in == 4) begin
					state<=4272;
					out<=83;
				end
			end
			2372: begin
				if(in == 0) begin
					state<=2373;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=6262;
					out<=86;
				end
				if(in == 3) begin
					state<=375;
					out<=87;
				end
				if(in == 4) begin
					state<=4273;
					out<=88;
				end
			end
			2373: begin
				if(in == 0) begin
					state<=2374;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=6263;
					out<=91;
				end
				if(in == 3) begin
					state<=376;
					out<=92;
				end
				if(in == 4) begin
					state<=4274;
					out<=93;
				end
			end
			2374: begin
				if(in == 0) begin
					state<=2375;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=6264;
					out<=96;
				end
				if(in == 3) begin
					state<=377;
					out<=97;
				end
				if(in == 4) begin
					state<=4275;
					out<=98;
				end
			end
			2375: begin
				if(in == 0) begin
					state<=2376;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=6265;
					out<=101;
				end
				if(in == 3) begin
					state<=378;
					out<=102;
				end
				if(in == 4) begin
					state<=4276;
					out<=103;
				end
			end
			2376: begin
				if(in == 0) begin
					state<=2377;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=6266;
					out<=106;
				end
				if(in == 3) begin
					state<=379;
					out<=107;
				end
				if(in == 4) begin
					state<=4277;
					out<=108;
				end
			end
			2377: begin
				if(in == 0) begin
					state<=2378;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=6267;
					out<=111;
				end
				if(in == 3) begin
					state<=380;
					out<=112;
				end
				if(in == 4) begin
					state<=4278;
					out<=113;
				end
			end
			2378: begin
				if(in == 0) begin
					state<=2379;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=6268;
					out<=116;
				end
				if(in == 3) begin
					state<=381;
					out<=117;
				end
				if(in == 4) begin
					state<=4279;
					out<=118;
				end
			end
			2379: begin
				if(in == 0) begin
					state<=2380;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=6269;
					out<=121;
				end
				if(in == 3) begin
					state<=382;
					out<=122;
				end
				if(in == 4) begin
					state<=4280;
					out<=123;
				end
			end
			2380: begin
				if(in == 0) begin
					state<=2381;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=6270;
					out<=126;
				end
				if(in == 3) begin
					state<=383;
					out<=127;
				end
				if(in == 4) begin
					state<=4281;
					out<=128;
				end
			end
			2381: begin
				if(in == 0) begin
					state<=2382;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=6271;
					out<=131;
				end
				if(in == 3) begin
					state<=384;
					out<=132;
				end
				if(in == 4) begin
					state<=4282;
					out<=133;
				end
			end
			2382: begin
				if(in == 0) begin
					state<=2383;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=6272;
					out<=136;
				end
				if(in == 3) begin
					state<=385;
					out<=137;
				end
				if(in == 4) begin
					state<=4283;
					out<=138;
				end
			end
			2383: begin
				if(in == 0) begin
					state<=2384;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=6273;
					out<=141;
				end
				if(in == 3) begin
					state<=386;
					out<=142;
				end
				if(in == 4) begin
					state<=4284;
					out<=143;
				end
			end
			2384: begin
				if(in == 0) begin
					state<=2385;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=6274;
					out<=146;
				end
				if(in == 3) begin
					state<=387;
					out<=147;
				end
				if(in == 4) begin
					state<=4285;
					out<=148;
				end
			end
			2385: begin
				if(in == 0) begin
					state<=2386;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=6275;
					out<=151;
				end
				if(in == 3) begin
					state<=388;
					out<=152;
				end
				if(in == 4) begin
					state<=4286;
					out<=153;
				end
			end
			2386: begin
				if(in == 0) begin
					state<=2387;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=6276;
					out<=156;
				end
				if(in == 3) begin
					state<=389;
					out<=157;
				end
				if(in == 4) begin
					state<=4287;
					out<=158;
				end
			end
			2387: begin
				if(in == 0) begin
					state<=2388;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=6277;
					out<=161;
				end
				if(in == 3) begin
					state<=390;
					out<=162;
				end
				if(in == 4) begin
					state<=4288;
					out<=163;
				end
			end
			2388: begin
				if(in == 0) begin
					state<=2389;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=6278;
					out<=166;
				end
				if(in == 3) begin
					state<=391;
					out<=167;
				end
				if(in == 4) begin
					state<=4289;
					out<=168;
				end
			end
			2389: begin
				if(in == 0) begin
					state<=2390;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=6279;
					out<=171;
				end
				if(in == 3) begin
					state<=392;
					out<=172;
				end
				if(in == 4) begin
					state<=4290;
					out<=173;
				end
			end
			2390: begin
				if(in == 0) begin
					state<=2391;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=6280;
					out<=176;
				end
				if(in == 3) begin
					state<=393;
					out<=177;
				end
				if(in == 4) begin
					state<=4291;
					out<=178;
				end
			end
			2391: begin
				if(in == 0) begin
					state<=2392;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=6281;
					out<=181;
				end
				if(in == 3) begin
					state<=394;
					out<=182;
				end
				if(in == 4) begin
					state<=4292;
					out<=183;
				end
			end
			2392: begin
				if(in == 0) begin
					state<=2393;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=6282;
					out<=186;
				end
				if(in == 3) begin
					state<=395;
					out<=187;
				end
				if(in == 4) begin
					state<=4293;
					out<=188;
				end
			end
			2393: begin
				if(in == 0) begin
					state<=3385;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=7274;
					out<=191;
				end
				if(in == 3) begin
					state<=999;
					out<=192;
				end
				if(in == 4) begin
					state<=4897;
					out<=193;
				end
			end
			2394: begin
				if(in == 0) begin
					state<=2395;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=6284;
					out<=196;
				end
				if(in == 3) begin
					state<=397;
					out<=197;
				end
				if(in == 4) begin
					state<=4295;
					out<=198;
				end
			end
			2395: begin
				if(in == 0) begin
					state<=2396;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=6285;
					out<=201;
				end
				if(in == 3) begin
					state<=398;
					out<=202;
				end
				if(in == 4) begin
					state<=4296;
					out<=203;
				end
			end
			2396: begin
				if(in == 0) begin
					state<=2397;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=6286;
					out<=206;
				end
				if(in == 3) begin
					state<=399;
					out<=207;
				end
				if(in == 4) begin
					state<=4297;
					out<=208;
				end
			end
			2397: begin
				if(in == 0) begin
					state<=2398;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=6287;
					out<=211;
				end
				if(in == 3) begin
					state<=400;
					out<=212;
				end
				if(in == 4) begin
					state<=4298;
					out<=213;
				end
			end
			2398: begin
				if(in == 0) begin
					state<=2399;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=6288;
					out<=216;
				end
				if(in == 3) begin
					state<=401;
					out<=217;
				end
				if(in == 4) begin
					state<=4299;
					out<=218;
				end
			end
			2399: begin
				if(in == 0) begin
					state<=2400;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=6289;
					out<=221;
				end
				if(in == 3) begin
					state<=402;
					out<=222;
				end
				if(in == 4) begin
					state<=4300;
					out<=223;
				end
			end
			2400: begin
				if(in == 0) begin
					state<=2401;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=6290;
					out<=226;
				end
				if(in == 3) begin
					state<=403;
					out<=227;
				end
				if(in == 4) begin
					state<=4301;
					out<=228;
				end
			end
			2401: begin
				if(in == 0) begin
					state<=2402;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=6291;
					out<=231;
				end
				if(in == 3) begin
					state<=404;
					out<=232;
				end
				if(in == 4) begin
					state<=4302;
					out<=233;
				end
			end
			2402: begin
				if(in == 0) begin
					state<=2403;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=6292;
					out<=236;
				end
				if(in == 3) begin
					state<=405;
					out<=237;
				end
				if(in == 4) begin
					state<=4303;
					out<=238;
				end
			end
			2403: begin
				if(in == 0) begin
					state<=2404;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=6293;
					out<=241;
				end
				if(in == 3) begin
					state<=406;
					out<=242;
				end
				if(in == 4) begin
					state<=4304;
					out<=243;
				end
			end
			2404: begin
				if(in == 0) begin
					state<=2405;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=6294;
					out<=246;
				end
				if(in == 3) begin
					state<=407;
					out<=247;
				end
				if(in == 4) begin
					state<=4305;
					out<=248;
				end
			end
			2405: begin
				if(in == 0) begin
					state<=2406;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=6295;
					out<=251;
				end
				if(in == 3) begin
					state<=408;
					out<=252;
				end
				if(in == 4) begin
					state<=4306;
					out<=253;
				end
			end
			2406: begin
				if(in == 0) begin
					state<=2407;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=6296;
					out<=0;
				end
				if(in == 3) begin
					state<=409;
					out<=1;
				end
				if(in == 4) begin
					state<=4307;
					out<=2;
				end
			end
			2407: begin
				if(in == 0) begin
					state<=2408;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=6297;
					out<=5;
				end
				if(in == 3) begin
					state<=410;
					out<=6;
				end
				if(in == 4) begin
					state<=4308;
					out<=7;
				end
			end
			2408: begin
				if(in == 0) begin
					state<=2409;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=6298;
					out<=10;
				end
				if(in == 3) begin
					state<=411;
					out<=11;
				end
				if(in == 4) begin
					state<=4309;
					out<=12;
				end
			end
			2409: begin
				if(in == 0) begin
					state<=2410;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=6299;
					out<=15;
				end
				if(in == 3) begin
					state<=412;
					out<=16;
				end
				if(in == 4) begin
					state<=4310;
					out<=17;
				end
			end
			2410: begin
				if(in == 0) begin
					state<=2411;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=6300;
					out<=20;
				end
				if(in == 3) begin
					state<=413;
					out<=21;
				end
				if(in == 4) begin
					state<=4311;
					out<=22;
				end
			end
			2411: begin
				if(in == 0) begin
					state<=2412;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=6301;
					out<=25;
				end
				if(in == 3) begin
					state<=414;
					out<=26;
				end
				if(in == 4) begin
					state<=4312;
					out<=27;
				end
			end
			2412: begin
				if(in == 0) begin
					state<=2413;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=6302;
					out<=30;
				end
				if(in == 3) begin
					state<=415;
					out<=31;
				end
				if(in == 4) begin
					state<=4313;
					out<=32;
				end
			end
			2413: begin
				if(in == 0) begin
					state<=2414;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=6303;
					out<=35;
				end
				if(in == 3) begin
					state<=416;
					out<=36;
				end
				if(in == 4) begin
					state<=4314;
					out<=37;
				end
			end
			2414: begin
				if(in == 0) begin
					state<=2415;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=6304;
					out<=40;
				end
				if(in == 3) begin
					state<=417;
					out<=41;
				end
				if(in == 4) begin
					state<=4315;
					out<=42;
				end
			end
			2415: begin
				if(in == 0) begin
					state<=2416;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=6305;
					out<=45;
				end
				if(in == 3) begin
					state<=418;
					out<=46;
				end
				if(in == 4) begin
					state<=4316;
					out<=47;
				end
			end
			2416: begin
				if(in == 0) begin
					state<=2417;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=6306;
					out<=50;
				end
				if(in == 3) begin
					state<=419;
					out<=51;
				end
				if(in == 4) begin
					state<=4317;
					out<=52;
				end
			end
			2417: begin
				if(in == 0) begin
					state<=2418;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=6307;
					out<=55;
				end
				if(in == 3) begin
					state<=420;
					out<=56;
				end
				if(in == 4) begin
					state<=4318;
					out<=57;
				end
			end
			2418: begin
				if(in == 0) begin
					state<=2419;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=6308;
					out<=60;
				end
				if(in == 3) begin
					state<=421;
					out<=61;
				end
				if(in == 4) begin
					state<=4319;
					out<=62;
				end
			end
			2419: begin
				if(in == 0) begin
					state<=2420;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=6309;
					out<=65;
				end
				if(in == 3) begin
					state<=422;
					out<=66;
				end
				if(in == 4) begin
					state<=4320;
					out<=67;
				end
			end
			2420: begin
				if(in == 0) begin
					state<=2421;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=6310;
					out<=70;
				end
				if(in == 3) begin
					state<=423;
					out<=71;
				end
				if(in == 4) begin
					state<=4321;
					out<=72;
				end
			end
			2421: begin
				if(in == 0) begin
					state<=2422;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=6311;
					out<=75;
				end
				if(in == 3) begin
					state<=424;
					out<=76;
				end
				if(in == 4) begin
					state<=4322;
					out<=77;
				end
			end
			2422: begin
				if(in == 0) begin
					state<=2423;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=6312;
					out<=80;
				end
				if(in == 3) begin
					state<=425;
					out<=81;
				end
				if(in == 4) begin
					state<=4323;
					out<=82;
				end
			end
			2423: begin
				if(in == 0) begin
					state<=2424;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=6313;
					out<=85;
				end
				if(in == 3) begin
					state<=426;
					out<=86;
				end
				if(in == 4) begin
					state<=4324;
					out<=87;
				end
			end
			2424: begin
				if(in == 0) begin
					state<=2425;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=6314;
					out<=90;
				end
				if(in == 3) begin
					state<=427;
					out<=91;
				end
				if(in == 4) begin
					state<=4325;
					out<=92;
				end
			end
			2425: begin
				if(in == 0) begin
					state<=2426;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=6315;
					out<=95;
				end
				if(in == 3) begin
					state<=428;
					out<=96;
				end
				if(in == 4) begin
					state<=4326;
					out<=97;
				end
			end
			2426: begin
				if(in == 0) begin
					state<=2427;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=6316;
					out<=100;
				end
				if(in == 3) begin
					state<=429;
					out<=101;
				end
				if(in == 4) begin
					state<=4327;
					out<=102;
				end
			end
			2427: begin
				if(in == 0) begin
					state<=2428;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=6317;
					out<=105;
				end
				if(in == 3) begin
					state<=430;
					out<=106;
				end
				if(in == 4) begin
					state<=4328;
					out<=107;
				end
			end
			2428: begin
				if(in == 0) begin
					state<=2429;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=6318;
					out<=110;
				end
				if(in == 3) begin
					state<=431;
					out<=111;
				end
				if(in == 4) begin
					state<=4329;
					out<=112;
				end
			end
			2429: begin
				if(in == 0) begin
					state<=2430;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=6319;
					out<=115;
				end
				if(in == 3) begin
					state<=432;
					out<=116;
				end
				if(in == 4) begin
					state<=4330;
					out<=117;
				end
			end
			2430: begin
				if(in == 0) begin
					state<=2431;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=6320;
					out<=120;
				end
				if(in == 3) begin
					state<=433;
					out<=121;
				end
				if(in == 4) begin
					state<=4331;
					out<=122;
				end
			end
			2431: begin
				if(in == 0) begin
					state<=2432;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=6321;
					out<=125;
				end
				if(in == 3) begin
					state<=434;
					out<=126;
				end
				if(in == 4) begin
					state<=4332;
					out<=127;
				end
			end
			2432: begin
				if(in == 0) begin
					state<=2433;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=6322;
					out<=130;
				end
				if(in == 3) begin
					state<=435;
					out<=131;
				end
				if(in == 4) begin
					state<=4333;
					out<=132;
				end
			end
			2433: begin
				if(in == 0) begin
					state<=2434;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=6323;
					out<=135;
				end
				if(in == 3) begin
					state<=436;
					out<=136;
				end
				if(in == 4) begin
					state<=4334;
					out<=137;
				end
			end
			2434: begin
				if(in == 0) begin
					state<=2435;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=6324;
					out<=140;
				end
				if(in == 3) begin
					state<=437;
					out<=141;
				end
				if(in == 4) begin
					state<=4335;
					out<=142;
				end
			end
			2435: begin
				if(in == 0) begin
					state<=2436;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=6325;
					out<=145;
				end
				if(in == 3) begin
					state<=438;
					out<=146;
				end
				if(in == 4) begin
					state<=4336;
					out<=147;
				end
			end
			2436: begin
				if(in == 0) begin
					state<=2437;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=6326;
					out<=150;
				end
				if(in == 3) begin
					state<=439;
					out<=151;
				end
				if(in == 4) begin
					state<=4337;
					out<=152;
				end
			end
			2437: begin
				if(in == 0) begin
					state<=2438;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=6327;
					out<=155;
				end
				if(in == 3) begin
					state<=440;
					out<=156;
				end
				if(in == 4) begin
					state<=4338;
					out<=157;
				end
			end
			2438: begin
				if(in == 0) begin
					state<=2439;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=6328;
					out<=160;
				end
				if(in == 3) begin
					state<=441;
					out<=161;
				end
				if(in == 4) begin
					state<=4339;
					out<=162;
				end
			end
			2439: begin
				if(in == 0) begin
					state<=2440;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=6329;
					out<=165;
				end
				if(in == 3) begin
					state<=442;
					out<=166;
				end
				if(in == 4) begin
					state<=4340;
					out<=167;
				end
			end
			2440: begin
				if(in == 0) begin
					state<=2441;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=6330;
					out<=170;
				end
				if(in == 3) begin
					state<=443;
					out<=171;
				end
				if(in == 4) begin
					state<=4341;
					out<=172;
				end
			end
			2441: begin
				if(in == 0) begin
					state<=2442;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=6331;
					out<=175;
				end
				if(in == 3) begin
					state<=444;
					out<=176;
				end
				if(in == 4) begin
					state<=4342;
					out<=177;
				end
			end
			2442: begin
				if(in == 0) begin
					state<=2443;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=6332;
					out<=180;
				end
				if(in == 3) begin
					state<=445;
					out<=181;
				end
				if(in == 4) begin
					state<=4343;
					out<=182;
				end
			end
			2443: begin
				if(in == 0) begin
					state<=2444;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=6333;
					out<=185;
				end
				if(in == 3) begin
					state<=446;
					out<=186;
				end
				if(in == 4) begin
					state<=4344;
					out<=187;
				end
			end
			2444: begin
				if(in == 0) begin
					state<=2445;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=6334;
					out<=190;
				end
				if(in == 3) begin
					state<=447;
					out<=191;
				end
				if(in == 4) begin
					state<=4345;
					out<=192;
				end
			end
			2445: begin
				if(in == 0) begin
					state<=2446;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=6335;
					out<=195;
				end
				if(in == 3) begin
					state<=448;
					out<=196;
				end
				if(in == 4) begin
					state<=4346;
					out<=197;
				end
			end
			2446: begin
				if(in == 0) begin
					state<=2447;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=6336;
					out<=200;
				end
				if(in == 3) begin
					state<=449;
					out<=201;
				end
				if(in == 4) begin
					state<=4347;
					out<=202;
				end
			end
			2447: begin
				if(in == 0) begin
					state<=2448;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=6337;
					out<=205;
				end
				if(in == 3) begin
					state<=450;
					out<=206;
				end
				if(in == 4) begin
					state<=4348;
					out<=207;
				end
			end
			2448: begin
				if(in == 0) begin
					state<=2449;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=6338;
					out<=210;
				end
				if(in == 3) begin
					state<=451;
					out<=211;
				end
				if(in == 4) begin
					state<=4349;
					out<=212;
				end
			end
			2449: begin
				if(in == 0) begin
					state<=2450;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=6339;
					out<=215;
				end
				if(in == 3) begin
					state<=452;
					out<=216;
				end
				if(in == 4) begin
					state<=4350;
					out<=217;
				end
			end
			2450: begin
				if(in == 0) begin
					state<=2451;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=6340;
					out<=220;
				end
				if(in == 3) begin
					state<=453;
					out<=221;
				end
				if(in == 4) begin
					state<=4351;
					out<=222;
				end
			end
			2451: begin
				if(in == 0) begin
					state<=2452;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=6341;
					out<=225;
				end
				if(in == 3) begin
					state<=454;
					out<=226;
				end
				if(in == 4) begin
					state<=4352;
					out<=227;
				end
			end
			2452: begin
				if(in == 0) begin
					state<=2453;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=6342;
					out<=230;
				end
				if(in == 3) begin
					state<=455;
					out<=231;
				end
				if(in == 4) begin
					state<=4353;
					out<=232;
				end
			end
			2453: begin
				if(in == 0) begin
					state<=2454;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=6343;
					out<=235;
				end
				if(in == 3) begin
					state<=456;
					out<=236;
				end
				if(in == 4) begin
					state<=4354;
					out<=237;
				end
			end
			2454: begin
				if(in == 0) begin
					state<=2455;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=6344;
					out<=240;
				end
				if(in == 3) begin
					state<=457;
					out<=241;
				end
				if(in == 4) begin
					state<=4355;
					out<=242;
				end
			end
			2455: begin
				if(in == 0) begin
					state<=2456;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=6345;
					out<=245;
				end
				if(in == 3) begin
					state<=458;
					out<=246;
				end
				if(in == 4) begin
					state<=4356;
					out<=247;
				end
			end
			2456: begin
				if(in == 0) begin
					state<=2457;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=6346;
					out<=250;
				end
				if(in == 3) begin
					state<=459;
					out<=251;
				end
				if(in == 4) begin
					state<=4357;
					out<=252;
				end
			end
			2457: begin
				if(in == 0) begin
					state<=2458;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=6347;
					out<=255;
				end
				if(in == 3) begin
					state<=460;
					out<=0;
				end
				if(in == 4) begin
					state<=4358;
					out<=1;
				end
			end
			2458: begin
				if(in == 0) begin
					state<=2459;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=6348;
					out<=4;
				end
				if(in == 3) begin
					state<=461;
					out<=5;
				end
				if(in == 4) begin
					state<=4359;
					out<=6;
				end
			end
			2459: begin
				if(in == 0) begin
					state<=2460;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=6349;
					out<=9;
				end
				if(in == 3) begin
					state<=462;
					out<=10;
				end
				if(in == 4) begin
					state<=4360;
					out<=11;
				end
			end
			2460: begin
				if(in == 0) begin
					state<=2461;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=6350;
					out<=14;
				end
				if(in == 3) begin
					state<=463;
					out<=15;
				end
				if(in == 4) begin
					state<=4361;
					out<=16;
				end
			end
			2461: begin
				if(in == 0) begin
					state<=2462;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=6351;
					out<=19;
				end
				if(in == 3) begin
					state<=464;
					out<=20;
				end
				if(in == 4) begin
					state<=4362;
					out<=21;
				end
			end
			2462: begin
				if(in == 0) begin
					state<=3416;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=7305;
					out<=24;
				end
				if(in == 3) begin
					state<=1484;
					out<=25;
				end
				if(in == 4) begin
					state<=5373;
					out<=26;
				end
			end
			2463: begin
				if(in == 0) begin
					state<=2464;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=6353;
					out<=29;
				end
				if(in == 3) begin
					state<=466;
					out<=30;
				end
				if(in == 4) begin
					state<=4364;
					out<=31;
				end
			end
			2464: begin
				if(in == 0) begin
					state<=2465;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=6354;
					out<=34;
				end
				if(in == 3) begin
					state<=467;
					out<=35;
				end
				if(in == 4) begin
					state<=4365;
					out<=36;
				end
			end
			2465: begin
				if(in == 0) begin
					state<=2466;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=6355;
					out<=39;
				end
				if(in == 3) begin
					state<=468;
					out<=40;
				end
				if(in == 4) begin
					state<=4366;
					out<=41;
				end
			end
			2466: begin
				if(in == 0) begin
					state<=2467;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=6356;
					out<=44;
				end
				if(in == 3) begin
					state<=469;
					out<=45;
				end
				if(in == 4) begin
					state<=4367;
					out<=46;
				end
			end
			2467: begin
				if(in == 0) begin
					state<=2468;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=6357;
					out<=49;
				end
				if(in == 3) begin
					state<=470;
					out<=50;
				end
				if(in == 4) begin
					state<=4368;
					out<=51;
				end
			end
			2468: begin
				if(in == 0) begin
					state<=2469;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=6358;
					out<=54;
				end
				if(in == 3) begin
					state<=471;
					out<=55;
				end
				if(in == 4) begin
					state<=4369;
					out<=56;
				end
			end
			2469: begin
				if(in == 0) begin
					state<=2470;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=6359;
					out<=59;
				end
				if(in == 3) begin
					state<=472;
					out<=60;
				end
				if(in == 4) begin
					state<=4370;
					out<=61;
				end
			end
			2470: begin
				if(in == 0) begin
					state<=2471;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=6360;
					out<=64;
				end
				if(in == 3) begin
					state<=473;
					out<=65;
				end
				if(in == 4) begin
					state<=4371;
					out<=66;
				end
			end
			2471: begin
				if(in == 0) begin
					state<=2472;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=6361;
					out<=69;
				end
				if(in == 3) begin
					state<=474;
					out<=70;
				end
				if(in == 4) begin
					state<=4372;
					out<=71;
				end
			end
			2472: begin
				if(in == 0) begin
					state<=2473;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=6362;
					out<=74;
				end
				if(in == 3) begin
					state<=475;
					out<=75;
				end
				if(in == 4) begin
					state<=4373;
					out<=76;
				end
			end
			2473: begin
				if(in == 0) begin
					state<=2474;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=6363;
					out<=79;
				end
				if(in == 3) begin
					state<=476;
					out<=80;
				end
				if(in == 4) begin
					state<=4374;
					out<=81;
				end
			end
			2474: begin
				if(in == 0) begin
					state<=2475;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=6364;
					out<=84;
				end
				if(in == 3) begin
					state<=477;
					out<=85;
				end
				if(in == 4) begin
					state<=4375;
					out<=86;
				end
			end
			2475: begin
				if(in == 0) begin
					state<=2476;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=6365;
					out<=89;
				end
				if(in == 3) begin
					state<=478;
					out<=90;
				end
				if(in == 4) begin
					state<=4376;
					out<=91;
				end
			end
			2476: begin
				if(in == 0) begin
					state<=2477;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=6366;
					out<=94;
				end
				if(in == 3) begin
					state<=479;
					out<=95;
				end
				if(in == 4) begin
					state<=4377;
					out<=96;
				end
			end
			2477: begin
				if(in == 0) begin
					state<=2478;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=6367;
					out<=99;
				end
				if(in == 3) begin
					state<=480;
					out<=100;
				end
				if(in == 4) begin
					state<=4378;
					out<=101;
				end
			end
			2478: begin
				if(in == 0) begin
					state<=2479;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=6368;
					out<=104;
				end
				if(in == 3) begin
					state<=481;
					out<=105;
				end
				if(in == 4) begin
					state<=4379;
					out<=106;
				end
			end
			2479: begin
				if(in == 0) begin
					state<=2480;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=6369;
					out<=109;
				end
				if(in == 3) begin
					state<=482;
					out<=110;
				end
				if(in == 4) begin
					state<=4380;
					out<=111;
				end
			end
			2480: begin
				if(in == 0) begin
					state<=2481;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=6370;
					out<=114;
				end
				if(in == 3) begin
					state<=483;
					out<=115;
				end
				if(in == 4) begin
					state<=4381;
					out<=116;
				end
			end
			2481: begin
				if(in == 0) begin
					state<=2482;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=6371;
					out<=119;
				end
				if(in == 3) begin
					state<=484;
					out<=120;
				end
				if(in == 4) begin
					state<=4382;
					out<=121;
				end
			end
			2482: begin
				if(in == 0) begin
					state<=2483;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=6372;
					out<=124;
				end
				if(in == 3) begin
					state<=485;
					out<=125;
				end
				if(in == 4) begin
					state<=4383;
					out<=126;
				end
			end
			2483: begin
				if(in == 0) begin
					state<=2484;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=6373;
					out<=129;
				end
				if(in == 3) begin
					state<=486;
					out<=130;
				end
				if(in == 4) begin
					state<=4384;
					out<=131;
				end
			end
			2484: begin
				if(in == 0) begin
					state<=2485;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=6374;
					out<=134;
				end
				if(in == 3) begin
					state<=487;
					out<=135;
				end
				if(in == 4) begin
					state<=4385;
					out<=136;
				end
			end
			2485: begin
				if(in == 0) begin
					state<=2486;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=6375;
					out<=139;
				end
				if(in == 3) begin
					state<=488;
					out<=140;
				end
				if(in == 4) begin
					state<=4386;
					out<=141;
				end
			end
			2486: begin
				if(in == 0) begin
					state<=2487;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=6376;
					out<=144;
				end
				if(in == 3) begin
					state<=489;
					out<=145;
				end
				if(in == 4) begin
					state<=4387;
					out<=146;
				end
			end
			2487: begin
				if(in == 0) begin
					state<=2488;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=6377;
					out<=149;
				end
				if(in == 3) begin
					state<=490;
					out<=150;
				end
				if(in == 4) begin
					state<=4388;
					out<=151;
				end
			end
			2488: begin
				if(in == 0) begin
					state<=2489;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=6378;
					out<=154;
				end
				if(in == 3) begin
					state<=491;
					out<=155;
				end
				if(in == 4) begin
					state<=4389;
					out<=156;
				end
			end
			2489: begin
				if(in == 0) begin
					state<=2490;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=6379;
					out<=159;
				end
				if(in == 3) begin
					state<=492;
					out<=160;
				end
				if(in == 4) begin
					state<=4390;
					out<=161;
				end
			end
			2490: begin
				if(in == 0) begin
					state<=2491;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=6380;
					out<=164;
				end
				if(in == 3) begin
					state<=493;
					out<=165;
				end
				if(in == 4) begin
					state<=4391;
					out<=166;
				end
			end
			2491: begin
				if(in == 0) begin
					state<=2492;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=6381;
					out<=169;
				end
				if(in == 3) begin
					state<=494;
					out<=170;
				end
				if(in == 4) begin
					state<=4392;
					out<=171;
				end
			end
			2492: begin
				if(in == 0) begin
					state<=2493;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=6382;
					out<=174;
				end
				if(in == 3) begin
					state<=495;
					out<=175;
				end
				if(in == 4) begin
					state<=4393;
					out<=176;
				end
			end
			2493: begin
				if(in == 0) begin
					state<=2494;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=6383;
					out<=179;
				end
				if(in == 3) begin
					state<=496;
					out<=180;
				end
				if(in == 4) begin
					state<=4394;
					out<=181;
				end
			end
			2494: begin
				if(in == 0) begin
					state<=2495;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=6384;
					out<=184;
				end
				if(in == 3) begin
					state<=497;
					out<=185;
				end
				if(in == 4) begin
					state<=4395;
					out<=186;
				end
			end
			2495: begin
				if(in == 0) begin
					state<=2496;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=6385;
					out<=189;
				end
				if(in == 3) begin
					state<=498;
					out<=190;
				end
				if(in == 4) begin
					state<=4396;
					out<=191;
				end
			end
			2496: begin
				if(in == 0) begin
					state<=2497;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=6386;
					out<=194;
				end
				if(in == 3) begin
					state<=499;
					out<=195;
				end
				if(in == 4) begin
					state<=4397;
					out<=196;
				end
			end
			2497: begin
				if(in == 0) begin
					state<=2498;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=6387;
					out<=199;
				end
				if(in == 3) begin
					state<=500;
					out<=200;
				end
				if(in == 4) begin
					state<=4398;
					out<=201;
				end
			end
			2498: begin
				if(in == 0) begin
					state<=2499;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=6388;
					out<=204;
				end
				if(in == 3) begin
					state<=501;
					out<=205;
				end
				if(in == 4) begin
					state<=4399;
					out<=206;
				end
			end
			2499: begin
				if(in == 0) begin
					state<=2500;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=6389;
					out<=209;
				end
				if(in == 3) begin
					state<=502;
					out<=210;
				end
				if(in == 4) begin
					state<=4400;
					out<=211;
				end
			end
			2500: begin
				if(in == 0) begin
					state<=2501;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=6390;
					out<=214;
				end
				if(in == 3) begin
					state<=503;
					out<=215;
				end
				if(in == 4) begin
					state<=4401;
					out<=216;
				end
			end
			2501: begin
				if(in == 0) begin
					state<=2502;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=6391;
					out<=219;
				end
				if(in == 3) begin
					state<=504;
					out<=220;
				end
				if(in == 4) begin
					state<=4402;
					out<=221;
				end
			end
			2502: begin
				if(in == 0) begin
					state<=2503;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=6392;
					out<=224;
				end
				if(in == 3) begin
					state<=505;
					out<=225;
				end
				if(in == 4) begin
					state<=4403;
					out<=226;
				end
			end
			2503: begin
				if(in == 0) begin
					state<=2504;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=6393;
					out<=229;
				end
				if(in == 3) begin
					state<=506;
					out<=230;
				end
				if(in == 4) begin
					state<=4404;
					out<=231;
				end
			end
			2504: begin
				if(in == 0) begin
					state<=2505;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=6394;
					out<=234;
				end
				if(in == 3) begin
					state<=507;
					out<=235;
				end
				if(in == 4) begin
					state<=4405;
					out<=236;
				end
			end
			2505: begin
				if(in == 0) begin
					state<=2506;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=6395;
					out<=239;
				end
				if(in == 3) begin
					state<=508;
					out<=240;
				end
				if(in == 4) begin
					state<=4406;
					out<=241;
				end
			end
			2506: begin
				if(in == 0) begin
					state<=2507;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=6396;
					out<=244;
				end
				if(in == 3) begin
					state<=509;
					out<=245;
				end
				if(in == 4) begin
					state<=4407;
					out<=246;
				end
			end
			2507: begin
				if(in == 0) begin
					state<=2508;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=6397;
					out<=249;
				end
				if(in == 3) begin
					state<=510;
					out<=250;
				end
				if(in == 4) begin
					state<=4408;
					out<=251;
				end
			end
			2508: begin
				if(in == 0) begin
					state<=2509;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=6398;
					out<=254;
				end
				if(in == 3) begin
					state<=511;
					out<=255;
				end
				if(in == 4) begin
					state<=4409;
					out<=0;
				end
			end
			2509: begin
				if(in == 0) begin
					state<=2510;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=6399;
					out<=3;
				end
				if(in == 3) begin
					state<=512;
					out<=4;
				end
				if(in == 4) begin
					state<=4410;
					out<=5;
				end
			end
			2510: begin
				if(in == 0) begin
					state<=2511;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=6400;
					out<=8;
				end
				if(in == 3) begin
					state<=513;
					out<=9;
				end
				if(in == 4) begin
					state<=4411;
					out<=10;
				end
			end
			2511: begin
				if(in == 0) begin
					state<=2512;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=6401;
					out<=13;
				end
				if(in == 3) begin
					state<=514;
					out<=14;
				end
				if(in == 4) begin
					state<=4412;
					out<=15;
				end
			end
			2512: begin
				if(in == 0) begin
					state<=2513;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=6402;
					out<=18;
				end
				if(in == 3) begin
					state<=515;
					out<=19;
				end
				if(in == 4) begin
					state<=4413;
					out<=20;
				end
			end
			2513: begin
				if(in == 0) begin
					state<=2514;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=6403;
					out<=23;
				end
				if(in == 3) begin
					state<=516;
					out<=24;
				end
				if(in == 4) begin
					state<=4414;
					out<=25;
				end
			end
			2514: begin
				if(in == 0) begin
					state<=2515;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=6404;
					out<=28;
				end
				if(in == 3) begin
					state<=517;
					out<=29;
				end
				if(in == 4) begin
					state<=4415;
					out<=30;
				end
			end
			2515: begin
				if(in == 0) begin
					state<=2516;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=6405;
					out<=33;
				end
				if(in == 3) begin
					state<=518;
					out<=34;
				end
				if(in == 4) begin
					state<=4416;
					out<=35;
				end
			end
			2516: begin
				if(in == 0) begin
					state<=2517;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=6406;
					out<=38;
				end
				if(in == 3) begin
					state<=519;
					out<=39;
				end
				if(in == 4) begin
					state<=4417;
					out<=40;
				end
			end
			2517: begin
				if(in == 0) begin
					state<=2518;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=6407;
					out<=43;
				end
				if(in == 3) begin
					state<=520;
					out<=44;
				end
				if(in == 4) begin
					state<=4418;
					out<=45;
				end
			end
			2518: begin
				if(in == 0) begin
					state<=2519;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=6408;
					out<=48;
				end
				if(in == 3) begin
					state<=521;
					out<=49;
				end
				if(in == 4) begin
					state<=4419;
					out<=50;
				end
			end
			2519: begin
				if(in == 0) begin
					state<=2520;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=6409;
					out<=53;
				end
				if(in == 3) begin
					state<=522;
					out<=54;
				end
				if(in == 4) begin
					state<=4420;
					out<=55;
				end
			end
			2520: begin
				if(in == 0) begin
					state<=2521;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=6410;
					out<=58;
				end
				if(in == 3) begin
					state<=523;
					out<=59;
				end
				if(in == 4) begin
					state<=4421;
					out<=60;
				end
			end
			2521: begin
				if(in == 0) begin
					state<=2522;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=6411;
					out<=63;
				end
				if(in == 3) begin
					state<=524;
					out<=64;
				end
				if(in == 4) begin
					state<=4422;
					out<=65;
				end
			end
			2522: begin
				if(in == 0) begin
					state<=2523;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=6412;
					out<=68;
				end
				if(in == 3) begin
					state<=525;
					out<=69;
				end
				if(in == 4) begin
					state<=4423;
					out<=70;
				end
			end
			2523: begin
				if(in == 0) begin
					state<=2524;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=6413;
					out<=73;
				end
				if(in == 3) begin
					state<=526;
					out<=74;
				end
				if(in == 4) begin
					state<=4424;
					out<=75;
				end
			end
			2524: begin
				if(in == 0) begin
					state<=2525;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=6414;
					out<=78;
				end
				if(in == 3) begin
					state<=527;
					out<=79;
				end
				if(in == 4) begin
					state<=4425;
					out<=80;
				end
			end
			2525: begin
				if(in == 0) begin
					state<=2526;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=6415;
					out<=83;
				end
				if(in == 3) begin
					state<=528;
					out<=84;
				end
				if(in == 4) begin
					state<=4426;
					out<=85;
				end
			end
			2526: begin
				if(in == 0) begin
					state<=2527;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=6416;
					out<=88;
				end
				if(in == 3) begin
					state<=529;
					out<=89;
				end
				if(in == 4) begin
					state<=4427;
					out<=90;
				end
			end
			2527: begin
				if(in == 0) begin
					state<=2528;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=6417;
					out<=93;
				end
				if(in == 3) begin
					state<=530;
					out<=94;
				end
				if(in == 4) begin
					state<=4428;
					out<=95;
				end
			end
			2528: begin
				if(in == 0) begin
					state<=2529;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=6418;
					out<=98;
				end
				if(in == 3) begin
					state<=531;
					out<=99;
				end
				if(in == 4) begin
					state<=4429;
					out<=100;
				end
			end
			2529: begin
				if(in == 0) begin
					state<=2530;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=6419;
					out<=103;
				end
				if(in == 3) begin
					state<=532;
					out<=104;
				end
				if(in == 4) begin
					state<=4430;
					out<=105;
				end
			end
			2530: begin
				if(in == 0) begin
					state<=2531;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=6420;
					out<=108;
				end
				if(in == 3) begin
					state<=533;
					out<=109;
				end
				if(in == 4) begin
					state<=4431;
					out<=110;
				end
			end
			2531: begin
				if(in == 0) begin
					state<=3447;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=7336;
					out<=113;
				end
				if(in == 3) begin
					state<=1515;
					out<=114;
				end
				if(in == 4) begin
					state<=5404;
					out<=115;
				end
			end
			2532: begin
				if(in == 0) begin
					state<=2533;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=6422;
					out<=118;
				end
				if(in == 3) begin
					state<=535;
					out<=119;
				end
				if(in == 4) begin
					state<=4433;
					out<=120;
				end
			end
			2533: begin
				if(in == 0) begin
					state<=2534;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=6423;
					out<=123;
				end
				if(in == 3) begin
					state<=536;
					out<=124;
				end
				if(in == 4) begin
					state<=4434;
					out<=125;
				end
			end
			2534: begin
				if(in == 0) begin
					state<=2535;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=6424;
					out<=128;
				end
				if(in == 3) begin
					state<=537;
					out<=129;
				end
				if(in == 4) begin
					state<=4435;
					out<=130;
				end
			end
			2535: begin
				if(in == 0) begin
					state<=2536;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=6425;
					out<=133;
				end
				if(in == 3) begin
					state<=538;
					out<=134;
				end
				if(in == 4) begin
					state<=4436;
					out<=135;
				end
			end
			2536: begin
				if(in == 0) begin
					state<=2537;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=6426;
					out<=138;
				end
				if(in == 3) begin
					state<=539;
					out<=139;
				end
				if(in == 4) begin
					state<=4437;
					out<=140;
				end
			end
			2537: begin
				if(in == 0) begin
					state<=2538;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=6427;
					out<=143;
				end
				if(in == 3) begin
					state<=540;
					out<=144;
				end
				if(in == 4) begin
					state<=4438;
					out<=145;
				end
			end
			2538: begin
				if(in == 0) begin
					state<=2539;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=6428;
					out<=148;
				end
				if(in == 3) begin
					state<=541;
					out<=149;
				end
				if(in == 4) begin
					state<=4439;
					out<=150;
				end
			end
			2539: begin
				if(in == 0) begin
					state<=2540;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=6429;
					out<=153;
				end
				if(in == 3) begin
					state<=542;
					out<=154;
				end
				if(in == 4) begin
					state<=4440;
					out<=155;
				end
			end
			2540: begin
				if(in == 0) begin
					state<=2541;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=6430;
					out<=158;
				end
				if(in == 3) begin
					state<=543;
					out<=159;
				end
				if(in == 4) begin
					state<=4441;
					out<=160;
				end
			end
			2541: begin
				if(in == 0) begin
					state<=2542;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=6431;
					out<=163;
				end
				if(in == 3) begin
					state<=544;
					out<=164;
				end
				if(in == 4) begin
					state<=4442;
					out<=165;
				end
			end
			2542: begin
				if(in == 0) begin
					state<=2543;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=6432;
					out<=168;
				end
				if(in == 3) begin
					state<=545;
					out<=169;
				end
				if(in == 4) begin
					state<=4443;
					out<=170;
				end
			end
			2543: begin
				if(in == 0) begin
					state<=2544;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=6433;
					out<=173;
				end
				if(in == 3) begin
					state<=546;
					out<=174;
				end
				if(in == 4) begin
					state<=4444;
					out<=175;
				end
			end
			2544: begin
				if(in == 0) begin
					state<=2545;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=6434;
					out<=178;
				end
				if(in == 3) begin
					state<=547;
					out<=179;
				end
				if(in == 4) begin
					state<=4445;
					out<=180;
				end
			end
			2545: begin
				if(in == 0) begin
					state<=2546;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=6435;
					out<=183;
				end
				if(in == 3) begin
					state<=548;
					out<=184;
				end
				if(in == 4) begin
					state<=4446;
					out<=185;
				end
			end
			2546: begin
				if(in == 0) begin
					state<=2547;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=6436;
					out<=188;
				end
				if(in == 3) begin
					state<=549;
					out<=189;
				end
				if(in == 4) begin
					state<=4447;
					out<=190;
				end
			end
			2547: begin
				if(in == 0) begin
					state<=2548;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=6437;
					out<=193;
				end
				if(in == 3) begin
					state<=550;
					out<=194;
				end
				if(in == 4) begin
					state<=4448;
					out<=195;
				end
			end
			2548: begin
				if(in == 0) begin
					state<=2549;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=6438;
					out<=198;
				end
				if(in == 3) begin
					state<=551;
					out<=199;
				end
				if(in == 4) begin
					state<=4449;
					out<=200;
				end
			end
			2549: begin
				if(in == 0) begin
					state<=2550;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=6439;
					out<=203;
				end
				if(in == 3) begin
					state<=552;
					out<=204;
				end
				if(in == 4) begin
					state<=4450;
					out<=205;
				end
			end
			2550: begin
				if(in == 0) begin
					state<=2551;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=6440;
					out<=208;
				end
				if(in == 3) begin
					state<=553;
					out<=209;
				end
				if(in == 4) begin
					state<=4451;
					out<=210;
				end
			end
			2551: begin
				if(in == 0) begin
					state<=2552;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=6441;
					out<=213;
				end
				if(in == 3) begin
					state<=554;
					out<=214;
				end
				if(in == 4) begin
					state<=4452;
					out<=215;
				end
			end
			2552: begin
				if(in == 0) begin
					state<=2553;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=6442;
					out<=218;
				end
				if(in == 3) begin
					state<=555;
					out<=219;
				end
				if(in == 4) begin
					state<=4453;
					out<=220;
				end
			end
			2553: begin
				if(in == 0) begin
					state<=2554;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=6443;
					out<=223;
				end
				if(in == 3) begin
					state<=556;
					out<=224;
				end
				if(in == 4) begin
					state<=4454;
					out<=225;
				end
			end
			2554: begin
				if(in == 0) begin
					state<=2555;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=6444;
					out<=228;
				end
				if(in == 3) begin
					state<=557;
					out<=229;
				end
				if(in == 4) begin
					state<=4455;
					out<=230;
				end
			end
			2555: begin
				if(in == 0) begin
					state<=2556;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=6445;
					out<=233;
				end
				if(in == 3) begin
					state<=558;
					out<=234;
				end
				if(in == 4) begin
					state<=4456;
					out<=235;
				end
			end
			2556: begin
				if(in == 0) begin
					state<=2557;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=6446;
					out<=238;
				end
				if(in == 3) begin
					state<=559;
					out<=239;
				end
				if(in == 4) begin
					state<=4457;
					out<=240;
				end
			end
			2557: begin
				if(in == 0) begin
					state<=2558;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=6447;
					out<=243;
				end
				if(in == 3) begin
					state<=560;
					out<=244;
				end
				if(in == 4) begin
					state<=4458;
					out<=245;
				end
			end
			2558: begin
				if(in == 0) begin
					state<=2559;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=6448;
					out<=248;
				end
				if(in == 3) begin
					state<=561;
					out<=249;
				end
				if(in == 4) begin
					state<=4459;
					out<=250;
				end
			end
			2559: begin
				if(in == 0) begin
					state<=2560;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=6449;
					out<=253;
				end
				if(in == 3) begin
					state<=562;
					out<=254;
				end
				if(in == 4) begin
					state<=4460;
					out<=255;
				end
			end
			2560: begin
				if(in == 0) begin
					state<=2561;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=6450;
					out<=2;
				end
				if(in == 3) begin
					state<=563;
					out<=3;
				end
				if(in == 4) begin
					state<=4461;
					out<=4;
				end
			end
			2561: begin
				if(in == 0) begin
					state<=2562;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=6451;
					out<=7;
				end
				if(in == 3) begin
					state<=564;
					out<=8;
				end
				if(in == 4) begin
					state<=4462;
					out<=9;
				end
			end
			2562: begin
				if(in == 0) begin
					state<=2563;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=6452;
					out<=12;
				end
				if(in == 3) begin
					state<=565;
					out<=13;
				end
				if(in == 4) begin
					state<=4463;
					out<=14;
				end
			end
			2563: begin
				if(in == 0) begin
					state<=2564;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=6453;
					out<=17;
				end
				if(in == 3) begin
					state<=566;
					out<=18;
				end
				if(in == 4) begin
					state<=4464;
					out<=19;
				end
			end
			2564: begin
				if(in == 0) begin
					state<=2565;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=6454;
					out<=22;
				end
				if(in == 3) begin
					state<=567;
					out<=23;
				end
				if(in == 4) begin
					state<=4465;
					out<=24;
				end
			end
			2565: begin
				if(in == 0) begin
					state<=2566;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=6455;
					out<=27;
				end
				if(in == 3) begin
					state<=568;
					out<=28;
				end
				if(in == 4) begin
					state<=4466;
					out<=29;
				end
			end
			2566: begin
				if(in == 0) begin
					state<=2567;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=6456;
					out<=32;
				end
				if(in == 3) begin
					state<=569;
					out<=33;
				end
				if(in == 4) begin
					state<=4467;
					out<=34;
				end
			end
			2567: begin
				if(in == 0) begin
					state<=2568;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=6457;
					out<=37;
				end
				if(in == 3) begin
					state<=570;
					out<=38;
				end
				if(in == 4) begin
					state<=4468;
					out<=39;
				end
			end
			2568: begin
				if(in == 0) begin
					state<=2569;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=6458;
					out<=42;
				end
				if(in == 3) begin
					state<=571;
					out<=43;
				end
				if(in == 4) begin
					state<=4469;
					out<=44;
				end
			end
			2569: begin
				if(in == 0) begin
					state<=2570;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=6459;
					out<=47;
				end
				if(in == 3) begin
					state<=572;
					out<=48;
				end
				if(in == 4) begin
					state<=4470;
					out<=49;
				end
			end
			2570: begin
				if(in == 0) begin
					state<=2571;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=6460;
					out<=52;
				end
				if(in == 3) begin
					state<=573;
					out<=53;
				end
				if(in == 4) begin
					state<=4471;
					out<=54;
				end
			end
			2571: begin
				if(in == 0) begin
					state<=2572;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=6461;
					out<=57;
				end
				if(in == 3) begin
					state<=574;
					out<=58;
				end
				if(in == 4) begin
					state<=4472;
					out<=59;
				end
			end
			2572: begin
				if(in == 0) begin
					state<=2573;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=6462;
					out<=62;
				end
				if(in == 3) begin
					state<=575;
					out<=63;
				end
				if(in == 4) begin
					state<=4473;
					out<=64;
				end
			end
			2573: begin
				if(in == 0) begin
					state<=2574;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=6463;
					out<=67;
				end
				if(in == 3) begin
					state<=576;
					out<=68;
				end
				if(in == 4) begin
					state<=4474;
					out<=69;
				end
			end
			2574: begin
				if(in == 0) begin
					state<=2575;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=6464;
					out<=72;
				end
				if(in == 3) begin
					state<=577;
					out<=73;
				end
				if(in == 4) begin
					state<=4475;
					out<=74;
				end
			end
			2575: begin
				if(in == 0) begin
					state<=2576;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=6465;
					out<=77;
				end
				if(in == 3) begin
					state<=578;
					out<=78;
				end
				if(in == 4) begin
					state<=4476;
					out<=79;
				end
			end
			2576: begin
				if(in == 0) begin
					state<=2577;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=6466;
					out<=82;
				end
				if(in == 3) begin
					state<=579;
					out<=83;
				end
				if(in == 4) begin
					state<=4477;
					out<=84;
				end
			end
			2577: begin
				if(in == 0) begin
					state<=2578;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=6467;
					out<=87;
				end
				if(in == 3) begin
					state<=580;
					out<=88;
				end
				if(in == 4) begin
					state<=4478;
					out<=89;
				end
			end
			2578: begin
				if(in == 0) begin
					state<=2579;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=6468;
					out<=92;
				end
				if(in == 3) begin
					state<=581;
					out<=93;
				end
				if(in == 4) begin
					state<=4479;
					out<=94;
				end
			end
			2579: begin
				if(in == 0) begin
					state<=2580;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=6469;
					out<=97;
				end
				if(in == 3) begin
					state<=582;
					out<=98;
				end
				if(in == 4) begin
					state<=4480;
					out<=99;
				end
			end
			2580: begin
				if(in == 0) begin
					state<=2581;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=6470;
					out<=102;
				end
				if(in == 3) begin
					state<=583;
					out<=103;
				end
				if(in == 4) begin
					state<=4481;
					out<=104;
				end
			end
			2581: begin
				if(in == 0) begin
					state<=2582;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=6471;
					out<=107;
				end
				if(in == 3) begin
					state<=584;
					out<=108;
				end
				if(in == 4) begin
					state<=4482;
					out<=109;
				end
			end
			2582: begin
				if(in == 0) begin
					state<=2583;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=6472;
					out<=112;
				end
				if(in == 3) begin
					state<=585;
					out<=113;
				end
				if(in == 4) begin
					state<=4483;
					out<=114;
				end
			end
			2583: begin
				if(in == 0) begin
					state<=2584;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=6473;
					out<=117;
				end
				if(in == 3) begin
					state<=586;
					out<=118;
				end
				if(in == 4) begin
					state<=4484;
					out<=119;
				end
			end
			2584: begin
				if(in == 0) begin
					state<=2585;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=6474;
					out<=122;
				end
				if(in == 3) begin
					state<=587;
					out<=123;
				end
				if(in == 4) begin
					state<=4485;
					out<=124;
				end
			end
			2585: begin
				if(in == 0) begin
					state<=2586;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=6475;
					out<=127;
				end
				if(in == 3) begin
					state<=588;
					out<=128;
				end
				if(in == 4) begin
					state<=4486;
					out<=129;
				end
			end
			2586: begin
				if(in == 0) begin
					state<=2587;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=6476;
					out<=132;
				end
				if(in == 3) begin
					state<=589;
					out<=133;
				end
				if(in == 4) begin
					state<=4487;
					out<=134;
				end
			end
			2587: begin
				if(in == 0) begin
					state<=2588;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=6477;
					out<=137;
				end
				if(in == 3) begin
					state<=590;
					out<=138;
				end
				if(in == 4) begin
					state<=4488;
					out<=139;
				end
			end
			2588: begin
				if(in == 0) begin
					state<=2589;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=6478;
					out<=142;
				end
				if(in == 3) begin
					state<=591;
					out<=143;
				end
				if(in == 4) begin
					state<=4489;
					out<=144;
				end
			end
			2589: begin
				if(in == 0) begin
					state<=2590;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=6479;
					out<=147;
				end
				if(in == 3) begin
					state<=592;
					out<=148;
				end
				if(in == 4) begin
					state<=4490;
					out<=149;
				end
			end
			2590: begin
				if(in == 0) begin
					state<=2591;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=6480;
					out<=152;
				end
				if(in == 3) begin
					state<=593;
					out<=153;
				end
				if(in == 4) begin
					state<=4491;
					out<=154;
				end
			end
			2591: begin
				if(in == 0) begin
					state<=2592;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=6481;
					out<=157;
				end
				if(in == 3) begin
					state<=594;
					out<=158;
				end
				if(in == 4) begin
					state<=4492;
					out<=159;
				end
			end
			2592: begin
				if(in == 0) begin
					state<=2593;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=6482;
					out<=162;
				end
				if(in == 3) begin
					state<=595;
					out<=163;
				end
				if(in == 4) begin
					state<=4493;
					out<=164;
				end
			end
			2593: begin
				if(in == 0) begin
					state<=2594;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=6483;
					out<=167;
				end
				if(in == 3) begin
					state<=596;
					out<=168;
				end
				if(in == 4) begin
					state<=4494;
					out<=169;
				end
			end
			2594: begin
				if(in == 0) begin
					state<=2595;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=6484;
					out<=172;
				end
				if(in == 3) begin
					state<=597;
					out<=173;
				end
				if(in == 4) begin
					state<=4495;
					out<=174;
				end
			end
			2595: begin
				if(in == 0) begin
					state<=2596;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=6485;
					out<=177;
				end
				if(in == 3) begin
					state<=598;
					out<=178;
				end
				if(in == 4) begin
					state<=4496;
					out<=179;
				end
			end
			2596: begin
				if(in == 0) begin
					state<=2597;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=6486;
					out<=182;
				end
				if(in == 3) begin
					state<=599;
					out<=183;
				end
				if(in == 4) begin
					state<=4497;
					out<=184;
				end
			end
			2597: begin
				if(in == 0) begin
					state<=2598;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=6487;
					out<=187;
				end
				if(in == 3) begin
					state<=600;
					out<=188;
				end
				if(in == 4) begin
					state<=4498;
					out<=189;
				end
			end
			2598: begin
				if(in == 0) begin
					state<=2599;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=6488;
					out<=192;
				end
				if(in == 3) begin
					state<=601;
					out<=193;
				end
				if(in == 4) begin
					state<=4499;
					out<=194;
				end
			end
			2599: begin
				if(in == 0) begin
					state<=2600;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=6489;
					out<=197;
				end
				if(in == 3) begin
					state<=602;
					out<=198;
				end
				if(in == 4) begin
					state<=4500;
					out<=199;
				end
			end
			2600: begin
				if(in == 0) begin
					state<=3478;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=7367;
					out<=202;
				end
				if(in == 3) begin
					state<=1546;
					out<=203;
				end
				if(in == 4) begin
					state<=5435;
					out<=204;
				end
			end
			2601: begin
				if(in == 0) begin
					state<=2602;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=6491;
					out<=207;
				end
				if(in == 3) begin
					state<=604;
					out<=208;
				end
				if(in == 4) begin
					state<=4502;
					out<=209;
				end
			end
			2602: begin
				if(in == 0) begin
					state<=2603;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=6492;
					out<=212;
				end
				if(in == 3) begin
					state<=605;
					out<=213;
				end
				if(in == 4) begin
					state<=4503;
					out<=214;
				end
			end
			2603: begin
				if(in == 0) begin
					state<=2604;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=6493;
					out<=217;
				end
				if(in == 3) begin
					state<=606;
					out<=218;
				end
				if(in == 4) begin
					state<=4504;
					out<=219;
				end
			end
			2604: begin
				if(in == 0) begin
					state<=2605;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=6494;
					out<=222;
				end
				if(in == 3) begin
					state<=607;
					out<=223;
				end
				if(in == 4) begin
					state<=4505;
					out<=224;
				end
			end
			2605: begin
				if(in == 0) begin
					state<=2606;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=6495;
					out<=227;
				end
				if(in == 3) begin
					state<=608;
					out<=228;
				end
				if(in == 4) begin
					state<=4506;
					out<=229;
				end
			end
			2606: begin
				if(in == 0) begin
					state<=2607;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=6496;
					out<=232;
				end
				if(in == 3) begin
					state<=609;
					out<=233;
				end
				if(in == 4) begin
					state<=4507;
					out<=234;
				end
			end
			2607: begin
				if(in == 0) begin
					state<=2608;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=6497;
					out<=237;
				end
				if(in == 3) begin
					state<=610;
					out<=238;
				end
				if(in == 4) begin
					state<=4508;
					out<=239;
				end
			end
			2608: begin
				if(in == 0) begin
					state<=2609;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=6498;
					out<=242;
				end
				if(in == 3) begin
					state<=611;
					out<=243;
				end
				if(in == 4) begin
					state<=4509;
					out<=244;
				end
			end
			2609: begin
				if(in == 0) begin
					state<=2610;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=6499;
					out<=247;
				end
				if(in == 3) begin
					state<=612;
					out<=248;
				end
				if(in == 4) begin
					state<=4510;
					out<=249;
				end
			end
			2610: begin
				if(in == 0) begin
					state<=2611;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=6500;
					out<=252;
				end
				if(in == 3) begin
					state<=613;
					out<=253;
				end
				if(in == 4) begin
					state<=4511;
					out<=254;
				end
			end
			2611: begin
				if(in == 0) begin
					state<=2612;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=6501;
					out<=1;
				end
				if(in == 3) begin
					state<=614;
					out<=2;
				end
				if(in == 4) begin
					state<=4512;
					out<=3;
				end
			end
			2612: begin
				if(in == 0) begin
					state<=2613;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=6502;
					out<=6;
				end
				if(in == 3) begin
					state<=615;
					out<=7;
				end
				if(in == 4) begin
					state<=4513;
					out<=8;
				end
			end
			2613: begin
				if(in == 0) begin
					state<=2614;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=6503;
					out<=11;
				end
				if(in == 3) begin
					state<=616;
					out<=12;
				end
				if(in == 4) begin
					state<=4514;
					out<=13;
				end
			end
			2614: begin
				if(in == 0) begin
					state<=2615;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=6504;
					out<=16;
				end
				if(in == 3) begin
					state<=617;
					out<=17;
				end
				if(in == 4) begin
					state<=4515;
					out<=18;
				end
			end
			2615: begin
				if(in == 0) begin
					state<=2616;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=6505;
					out<=21;
				end
				if(in == 3) begin
					state<=618;
					out<=22;
				end
				if(in == 4) begin
					state<=4516;
					out<=23;
				end
			end
			2616: begin
				if(in == 0) begin
					state<=2617;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=6506;
					out<=26;
				end
				if(in == 3) begin
					state<=619;
					out<=27;
				end
				if(in == 4) begin
					state<=4517;
					out<=28;
				end
			end
			2617: begin
				if(in == 0) begin
					state<=2618;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=6507;
					out<=31;
				end
				if(in == 3) begin
					state<=620;
					out<=32;
				end
				if(in == 4) begin
					state<=4518;
					out<=33;
				end
			end
			2618: begin
				if(in == 0) begin
					state<=2619;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=6508;
					out<=36;
				end
				if(in == 3) begin
					state<=621;
					out<=37;
				end
				if(in == 4) begin
					state<=4519;
					out<=38;
				end
			end
			2619: begin
				if(in == 0) begin
					state<=2620;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=6509;
					out<=41;
				end
				if(in == 3) begin
					state<=622;
					out<=42;
				end
				if(in == 4) begin
					state<=4520;
					out<=43;
				end
			end
			2620: begin
				if(in == 0) begin
					state<=2621;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=6510;
					out<=46;
				end
				if(in == 3) begin
					state<=623;
					out<=47;
				end
				if(in == 4) begin
					state<=4521;
					out<=48;
				end
			end
			2621: begin
				if(in == 0) begin
					state<=2622;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=6511;
					out<=51;
				end
				if(in == 3) begin
					state<=624;
					out<=52;
				end
				if(in == 4) begin
					state<=4522;
					out<=53;
				end
			end
			2622: begin
				if(in == 0) begin
					state<=2623;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=6512;
					out<=56;
				end
				if(in == 3) begin
					state<=625;
					out<=57;
				end
				if(in == 4) begin
					state<=4523;
					out<=58;
				end
			end
			2623: begin
				if(in == 0) begin
					state<=2624;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=6513;
					out<=61;
				end
				if(in == 3) begin
					state<=626;
					out<=62;
				end
				if(in == 4) begin
					state<=4524;
					out<=63;
				end
			end
			2624: begin
				if(in == 0) begin
					state<=2625;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=6514;
					out<=66;
				end
				if(in == 3) begin
					state<=627;
					out<=67;
				end
				if(in == 4) begin
					state<=4525;
					out<=68;
				end
			end
			2625: begin
				if(in == 0) begin
					state<=2626;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=6515;
					out<=71;
				end
				if(in == 3) begin
					state<=628;
					out<=72;
				end
				if(in == 4) begin
					state<=4526;
					out<=73;
				end
			end
			2626: begin
				if(in == 0) begin
					state<=2627;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=6516;
					out<=76;
				end
				if(in == 3) begin
					state<=629;
					out<=77;
				end
				if(in == 4) begin
					state<=4527;
					out<=78;
				end
			end
			2627: begin
				if(in == 0) begin
					state<=2628;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=6517;
					out<=81;
				end
				if(in == 3) begin
					state<=630;
					out<=82;
				end
				if(in == 4) begin
					state<=4528;
					out<=83;
				end
			end
			2628: begin
				if(in == 0) begin
					state<=2629;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=6518;
					out<=86;
				end
				if(in == 3) begin
					state<=631;
					out<=87;
				end
				if(in == 4) begin
					state<=4529;
					out<=88;
				end
			end
			2629: begin
				if(in == 0) begin
					state<=2630;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=6519;
					out<=91;
				end
				if(in == 3) begin
					state<=632;
					out<=92;
				end
				if(in == 4) begin
					state<=4530;
					out<=93;
				end
			end
			2630: begin
				if(in == 0) begin
					state<=2631;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=6520;
					out<=96;
				end
				if(in == 3) begin
					state<=633;
					out<=97;
				end
				if(in == 4) begin
					state<=4531;
					out<=98;
				end
			end
			2631: begin
				if(in == 0) begin
					state<=2632;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=6521;
					out<=101;
				end
				if(in == 3) begin
					state<=634;
					out<=102;
				end
				if(in == 4) begin
					state<=4532;
					out<=103;
				end
			end
			2632: begin
				if(in == 0) begin
					state<=2633;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=6522;
					out<=106;
				end
				if(in == 3) begin
					state<=635;
					out<=107;
				end
				if(in == 4) begin
					state<=4533;
					out<=108;
				end
			end
			2633: begin
				if(in == 0) begin
					state<=2634;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=6523;
					out<=111;
				end
				if(in == 3) begin
					state<=636;
					out<=112;
				end
				if(in == 4) begin
					state<=4534;
					out<=113;
				end
			end
			2634: begin
				if(in == 0) begin
					state<=2635;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=6524;
					out<=116;
				end
				if(in == 3) begin
					state<=637;
					out<=117;
				end
				if(in == 4) begin
					state<=4535;
					out<=118;
				end
			end
			2635: begin
				if(in == 0) begin
					state<=2636;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=6525;
					out<=121;
				end
				if(in == 3) begin
					state<=638;
					out<=122;
				end
				if(in == 4) begin
					state<=4536;
					out<=123;
				end
			end
			2636: begin
				if(in == 0) begin
					state<=2637;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=6526;
					out<=126;
				end
				if(in == 3) begin
					state<=639;
					out<=127;
				end
				if(in == 4) begin
					state<=4537;
					out<=128;
				end
			end
			2637: begin
				if(in == 0) begin
					state<=2638;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=6527;
					out<=131;
				end
				if(in == 3) begin
					state<=640;
					out<=132;
				end
				if(in == 4) begin
					state<=4538;
					out<=133;
				end
			end
			2638: begin
				if(in == 0) begin
					state<=2639;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=6528;
					out<=136;
				end
				if(in == 3) begin
					state<=641;
					out<=137;
				end
				if(in == 4) begin
					state<=4539;
					out<=138;
				end
			end
			2639: begin
				if(in == 0) begin
					state<=2640;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=6529;
					out<=141;
				end
				if(in == 3) begin
					state<=642;
					out<=142;
				end
				if(in == 4) begin
					state<=4540;
					out<=143;
				end
			end
			2640: begin
				if(in == 0) begin
					state<=2641;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=6530;
					out<=146;
				end
				if(in == 3) begin
					state<=643;
					out<=147;
				end
				if(in == 4) begin
					state<=4541;
					out<=148;
				end
			end
			2641: begin
				if(in == 0) begin
					state<=2642;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=6531;
					out<=151;
				end
				if(in == 3) begin
					state<=644;
					out<=152;
				end
				if(in == 4) begin
					state<=4542;
					out<=153;
				end
			end
			2642: begin
				if(in == 0) begin
					state<=2643;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=6532;
					out<=156;
				end
				if(in == 3) begin
					state<=645;
					out<=157;
				end
				if(in == 4) begin
					state<=4543;
					out<=158;
				end
			end
			2643: begin
				if(in == 0) begin
					state<=2644;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=6533;
					out<=161;
				end
				if(in == 3) begin
					state<=646;
					out<=162;
				end
				if(in == 4) begin
					state<=4544;
					out<=163;
				end
			end
			2644: begin
				if(in == 0) begin
					state<=2645;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=6534;
					out<=166;
				end
				if(in == 3) begin
					state<=647;
					out<=167;
				end
				if(in == 4) begin
					state<=4545;
					out<=168;
				end
			end
			2645: begin
				if(in == 0) begin
					state<=2646;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=6535;
					out<=171;
				end
				if(in == 3) begin
					state<=648;
					out<=172;
				end
				if(in == 4) begin
					state<=4546;
					out<=173;
				end
			end
			2646: begin
				if(in == 0) begin
					state<=2647;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=6536;
					out<=176;
				end
				if(in == 3) begin
					state<=649;
					out<=177;
				end
				if(in == 4) begin
					state<=4547;
					out<=178;
				end
			end
			2647: begin
				if(in == 0) begin
					state<=2648;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=6537;
					out<=181;
				end
				if(in == 3) begin
					state<=650;
					out<=182;
				end
				if(in == 4) begin
					state<=4548;
					out<=183;
				end
			end
			2648: begin
				if(in == 0) begin
					state<=2649;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=6538;
					out<=186;
				end
				if(in == 3) begin
					state<=651;
					out<=187;
				end
				if(in == 4) begin
					state<=4549;
					out<=188;
				end
			end
			2649: begin
				if(in == 0) begin
					state<=2650;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=6539;
					out<=191;
				end
				if(in == 3) begin
					state<=652;
					out<=192;
				end
				if(in == 4) begin
					state<=4550;
					out<=193;
				end
			end
			2650: begin
				if(in == 0) begin
					state<=2651;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=6540;
					out<=196;
				end
				if(in == 3) begin
					state<=653;
					out<=197;
				end
				if(in == 4) begin
					state<=4551;
					out<=198;
				end
			end
			2651: begin
				if(in == 0) begin
					state<=2652;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=6541;
					out<=201;
				end
				if(in == 3) begin
					state<=654;
					out<=202;
				end
				if(in == 4) begin
					state<=4552;
					out<=203;
				end
			end
			2652: begin
				if(in == 0) begin
					state<=2653;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=6542;
					out<=206;
				end
				if(in == 3) begin
					state<=655;
					out<=207;
				end
				if(in == 4) begin
					state<=4553;
					out<=208;
				end
			end
			2653: begin
				if(in == 0) begin
					state<=2654;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=6543;
					out<=211;
				end
				if(in == 3) begin
					state<=656;
					out<=212;
				end
				if(in == 4) begin
					state<=4554;
					out<=213;
				end
			end
			2654: begin
				if(in == 0) begin
					state<=2655;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=6544;
					out<=216;
				end
				if(in == 3) begin
					state<=657;
					out<=217;
				end
				if(in == 4) begin
					state<=4555;
					out<=218;
				end
			end
			2655: begin
				if(in == 0) begin
					state<=2656;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=6545;
					out<=221;
				end
				if(in == 3) begin
					state<=658;
					out<=222;
				end
				if(in == 4) begin
					state<=4556;
					out<=223;
				end
			end
			2656: begin
				if(in == 0) begin
					state<=2657;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=6546;
					out<=226;
				end
				if(in == 3) begin
					state<=659;
					out<=227;
				end
				if(in == 4) begin
					state<=4557;
					out<=228;
				end
			end
			2657: begin
				if(in == 0) begin
					state<=2658;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=6547;
					out<=231;
				end
				if(in == 3) begin
					state<=660;
					out<=232;
				end
				if(in == 4) begin
					state<=4558;
					out<=233;
				end
			end
			2658: begin
				if(in == 0) begin
					state<=2659;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=6548;
					out<=236;
				end
				if(in == 3) begin
					state<=661;
					out<=237;
				end
				if(in == 4) begin
					state<=4559;
					out<=238;
				end
			end
			2659: begin
				if(in == 0) begin
					state<=2660;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=6549;
					out<=241;
				end
				if(in == 3) begin
					state<=662;
					out<=242;
				end
				if(in == 4) begin
					state<=4560;
					out<=243;
				end
			end
			2660: begin
				if(in == 0) begin
					state<=2661;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=6550;
					out<=246;
				end
				if(in == 3) begin
					state<=663;
					out<=247;
				end
				if(in == 4) begin
					state<=4561;
					out<=248;
				end
			end
			2661: begin
				if(in == 0) begin
					state<=2662;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=6551;
					out<=251;
				end
				if(in == 3) begin
					state<=664;
					out<=252;
				end
				if(in == 4) begin
					state<=4562;
					out<=253;
				end
			end
			2662: begin
				if(in == 0) begin
					state<=2663;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=6552;
					out<=0;
				end
				if(in == 3) begin
					state<=665;
					out<=1;
				end
				if(in == 4) begin
					state<=4563;
					out<=2;
				end
			end
			2663: begin
				if(in == 0) begin
					state<=2664;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=6553;
					out<=5;
				end
				if(in == 3) begin
					state<=666;
					out<=6;
				end
				if(in == 4) begin
					state<=4564;
					out<=7;
				end
			end
			2664: begin
				if(in == 0) begin
					state<=2665;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=6554;
					out<=10;
				end
				if(in == 3) begin
					state<=667;
					out<=11;
				end
				if(in == 4) begin
					state<=4565;
					out<=12;
				end
			end
			2665: begin
				if(in == 0) begin
					state<=2666;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=6555;
					out<=15;
				end
				if(in == 3) begin
					state<=668;
					out<=16;
				end
				if(in == 4) begin
					state<=4566;
					out<=17;
				end
			end
			2666: begin
				if(in == 0) begin
					state<=2667;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=6556;
					out<=20;
				end
				if(in == 3) begin
					state<=669;
					out<=21;
				end
				if(in == 4) begin
					state<=4567;
					out<=22;
				end
			end
			2667: begin
				if(in == 0) begin
					state<=2668;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=6557;
					out<=25;
				end
				if(in == 3) begin
					state<=670;
					out<=26;
				end
				if(in == 4) begin
					state<=4568;
					out<=27;
				end
			end
			2668: begin
				if(in == 0) begin
					state<=2669;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=6558;
					out<=30;
				end
				if(in == 3) begin
					state<=671;
					out<=31;
				end
				if(in == 4) begin
					state<=4569;
					out<=32;
				end
			end
			2669: begin
				if(in == 0) begin
					state<=3230;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=7119;
					out<=35;
				end
				if(in == 3) begin
					state<=1577;
					out<=36;
				end
				if(in == 4) begin
					state<=5466;
					out<=37;
				end
			end
			2670: begin
				if(in == 0) begin
					state<=2671;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=6560;
					out<=40;
				end
				if(in == 3) begin
					state<=673;
					out<=41;
				end
				if(in == 4) begin
					state<=4571;
					out<=42;
				end
			end
			2671: begin
				if(in == 0) begin
					state<=2672;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=6561;
					out<=45;
				end
				if(in == 3) begin
					state<=674;
					out<=46;
				end
				if(in == 4) begin
					state<=4572;
					out<=47;
				end
			end
			2672: begin
				if(in == 0) begin
					state<=2673;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=6562;
					out<=50;
				end
				if(in == 3) begin
					state<=675;
					out<=51;
				end
				if(in == 4) begin
					state<=4573;
					out<=52;
				end
			end
			2673: begin
				if(in == 0) begin
					state<=2674;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=6563;
					out<=55;
				end
				if(in == 3) begin
					state<=676;
					out<=56;
				end
				if(in == 4) begin
					state<=4574;
					out<=57;
				end
			end
			2674: begin
				if(in == 0) begin
					state<=2675;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=6564;
					out<=60;
				end
				if(in == 3) begin
					state<=677;
					out<=61;
				end
				if(in == 4) begin
					state<=4575;
					out<=62;
				end
			end
			2675: begin
				if(in == 0) begin
					state<=2676;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=6565;
					out<=65;
				end
				if(in == 3) begin
					state<=678;
					out<=66;
				end
				if(in == 4) begin
					state<=4576;
					out<=67;
				end
			end
			2676: begin
				if(in == 0) begin
					state<=2677;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=6566;
					out<=70;
				end
				if(in == 3) begin
					state<=679;
					out<=71;
				end
				if(in == 4) begin
					state<=4577;
					out<=72;
				end
			end
			2677: begin
				if(in == 0) begin
					state<=2678;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=6567;
					out<=75;
				end
				if(in == 3) begin
					state<=680;
					out<=76;
				end
				if(in == 4) begin
					state<=4578;
					out<=77;
				end
			end
			2678: begin
				if(in == 0) begin
					state<=2679;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=6568;
					out<=80;
				end
				if(in == 3) begin
					state<=681;
					out<=81;
				end
				if(in == 4) begin
					state<=4579;
					out<=82;
				end
			end
			2679: begin
				if(in == 0) begin
					state<=2680;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=6569;
					out<=85;
				end
				if(in == 3) begin
					state<=682;
					out<=86;
				end
				if(in == 4) begin
					state<=4580;
					out<=87;
				end
			end
			2680: begin
				if(in == 0) begin
					state<=2681;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=6570;
					out<=90;
				end
				if(in == 3) begin
					state<=683;
					out<=91;
				end
				if(in == 4) begin
					state<=4581;
					out<=92;
				end
			end
			2681: begin
				if(in == 0) begin
					state<=2682;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=6571;
					out<=95;
				end
				if(in == 3) begin
					state<=684;
					out<=96;
				end
				if(in == 4) begin
					state<=4582;
					out<=97;
				end
			end
			2682: begin
				if(in == 0) begin
					state<=2683;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=6572;
					out<=100;
				end
				if(in == 3) begin
					state<=685;
					out<=101;
				end
				if(in == 4) begin
					state<=4583;
					out<=102;
				end
			end
			2683: begin
				if(in == 0) begin
					state<=2684;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=6573;
					out<=105;
				end
				if(in == 3) begin
					state<=686;
					out<=106;
				end
				if(in == 4) begin
					state<=4584;
					out<=107;
				end
			end
			2684: begin
				if(in == 0) begin
					state<=2685;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=6574;
					out<=110;
				end
				if(in == 3) begin
					state<=687;
					out<=111;
				end
				if(in == 4) begin
					state<=4585;
					out<=112;
				end
			end
			2685: begin
				if(in == 0) begin
					state<=2686;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=6575;
					out<=115;
				end
				if(in == 3) begin
					state<=688;
					out<=116;
				end
				if(in == 4) begin
					state<=4586;
					out<=117;
				end
			end
			2686: begin
				if(in == 0) begin
					state<=2687;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=6576;
					out<=120;
				end
				if(in == 3) begin
					state<=689;
					out<=121;
				end
				if(in == 4) begin
					state<=4587;
					out<=122;
				end
			end
			2687: begin
				if(in == 0) begin
					state<=2688;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=6577;
					out<=125;
				end
				if(in == 3) begin
					state<=690;
					out<=126;
				end
				if(in == 4) begin
					state<=4588;
					out<=127;
				end
			end
			2688: begin
				if(in == 0) begin
					state<=1999;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=5888;
					out<=130;
				end
				if(in == 3) begin
					state<=1;
					out<=131;
				end
				if(in == 4) begin
					state<=3899;
					out<=132;
				end
			end
			2689: begin
				if(in == 0) begin
					state<=2690;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=6579;
					out<=135;
				end
				if(in == 3) begin
					state<=692;
					out<=136;
				end
				if(in == 4) begin
					state<=4590;
					out<=137;
				end
			end
			2690: begin
				if(in == 0) begin
					state<=2691;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=6580;
					out<=140;
				end
				if(in == 3) begin
					state<=693;
					out<=141;
				end
				if(in == 4) begin
					state<=4591;
					out<=142;
				end
			end
			2691: begin
				if(in == 0) begin
					state<=2692;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=6581;
					out<=145;
				end
				if(in == 3) begin
					state<=694;
					out<=146;
				end
				if(in == 4) begin
					state<=4592;
					out<=147;
				end
			end
			2692: begin
				if(in == 0) begin
					state<=2693;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=6582;
					out<=150;
				end
				if(in == 3) begin
					state<=695;
					out<=151;
				end
				if(in == 4) begin
					state<=4593;
					out<=152;
				end
			end
			2693: begin
				if(in == 0) begin
					state<=2694;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=6583;
					out<=155;
				end
				if(in == 3) begin
					state<=696;
					out<=156;
				end
				if(in == 4) begin
					state<=4594;
					out<=157;
				end
			end
			2694: begin
				if(in == 0) begin
					state<=2695;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=6584;
					out<=160;
				end
				if(in == 3) begin
					state<=697;
					out<=161;
				end
				if(in == 4) begin
					state<=4595;
					out<=162;
				end
			end
			2695: begin
				if(in == 0) begin
					state<=2696;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=6585;
					out<=165;
				end
				if(in == 3) begin
					state<=698;
					out<=166;
				end
				if(in == 4) begin
					state<=4596;
					out<=167;
				end
			end
			2696: begin
				if(in == 0) begin
					state<=2697;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=6586;
					out<=170;
				end
				if(in == 3) begin
					state<=699;
					out<=171;
				end
				if(in == 4) begin
					state<=4597;
					out<=172;
				end
			end
			2697: begin
				if(in == 0) begin
					state<=2698;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=6587;
					out<=175;
				end
				if(in == 3) begin
					state<=700;
					out<=176;
				end
				if(in == 4) begin
					state<=4598;
					out<=177;
				end
			end
			2698: begin
				if(in == 0) begin
					state<=2699;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=6588;
					out<=180;
				end
				if(in == 3) begin
					state<=701;
					out<=181;
				end
				if(in == 4) begin
					state<=4599;
					out<=182;
				end
			end
			2699: begin
				if(in == 0) begin
					state<=2700;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=6589;
					out<=185;
				end
				if(in == 3) begin
					state<=702;
					out<=186;
				end
				if(in == 4) begin
					state<=4600;
					out<=187;
				end
			end
			2700: begin
				if(in == 0) begin
					state<=2701;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=6590;
					out<=190;
				end
				if(in == 3) begin
					state<=703;
					out<=191;
				end
				if(in == 4) begin
					state<=4601;
					out<=192;
				end
			end
			2701: begin
				if(in == 0) begin
					state<=2702;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=6591;
					out<=195;
				end
				if(in == 3) begin
					state<=704;
					out<=196;
				end
				if(in == 4) begin
					state<=4602;
					out<=197;
				end
			end
			2702: begin
				if(in == 0) begin
					state<=2703;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=6592;
					out<=200;
				end
				if(in == 3) begin
					state<=705;
					out<=201;
				end
				if(in == 4) begin
					state<=4603;
					out<=202;
				end
			end
			2703: begin
				if(in == 0) begin
					state<=2704;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=6593;
					out<=205;
				end
				if(in == 3) begin
					state<=706;
					out<=206;
				end
				if(in == 4) begin
					state<=4604;
					out<=207;
				end
			end
			2704: begin
				if(in == 0) begin
					state<=2705;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=6594;
					out<=210;
				end
				if(in == 3) begin
					state<=707;
					out<=211;
				end
				if(in == 4) begin
					state<=4605;
					out<=212;
				end
			end
			2705: begin
				if(in == 0) begin
					state<=2706;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=6595;
					out<=215;
				end
				if(in == 3) begin
					state<=708;
					out<=216;
				end
				if(in == 4) begin
					state<=4606;
					out<=217;
				end
			end
			2706: begin
				if(in == 0) begin
					state<=2707;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=6596;
					out<=220;
				end
				if(in == 3) begin
					state<=709;
					out<=221;
				end
				if(in == 4) begin
					state<=4607;
					out<=222;
				end
			end
			2707: begin
				if(in == 0) begin
					state<=2708;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=6597;
					out<=225;
				end
				if(in == 3) begin
					state<=710;
					out<=226;
				end
				if(in == 4) begin
					state<=4608;
					out<=227;
				end
			end
			2708: begin
				if(in == 0) begin
					state<=2709;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=6598;
					out<=230;
				end
				if(in == 3) begin
					state<=711;
					out<=231;
				end
				if(in == 4) begin
					state<=4609;
					out<=232;
				end
			end
			2709: begin
				if(in == 0) begin
					state<=2710;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=6599;
					out<=235;
				end
				if(in == 3) begin
					state<=712;
					out<=236;
				end
				if(in == 4) begin
					state<=4610;
					out<=237;
				end
			end
			2710: begin
				if(in == 0) begin
					state<=2711;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=6600;
					out<=240;
				end
				if(in == 3) begin
					state<=713;
					out<=241;
				end
				if(in == 4) begin
					state<=4611;
					out<=242;
				end
			end
			2711: begin
				if(in == 0) begin
					state<=2712;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=6601;
					out<=245;
				end
				if(in == 3) begin
					state<=714;
					out<=246;
				end
				if(in == 4) begin
					state<=4612;
					out<=247;
				end
			end
			2712: begin
				if(in == 0) begin
					state<=2713;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=6602;
					out<=250;
				end
				if(in == 3) begin
					state<=715;
					out<=251;
				end
				if(in == 4) begin
					state<=4613;
					out<=252;
				end
			end
			2713: begin
				if(in == 0) begin
					state<=2714;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=6603;
					out<=255;
				end
				if(in == 3) begin
					state<=716;
					out<=0;
				end
				if(in == 4) begin
					state<=4614;
					out<=1;
				end
			end
			2714: begin
				if(in == 0) begin
					state<=2715;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=6604;
					out<=4;
				end
				if(in == 3) begin
					state<=717;
					out<=5;
				end
				if(in == 4) begin
					state<=4615;
					out<=6;
				end
			end
			2715: begin
				if(in == 0) begin
					state<=2716;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=6605;
					out<=9;
				end
				if(in == 3) begin
					state<=718;
					out<=10;
				end
				if(in == 4) begin
					state<=4616;
					out<=11;
				end
			end
			2716: begin
				if(in == 0) begin
					state<=2717;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=6606;
					out<=14;
				end
				if(in == 3) begin
					state<=719;
					out<=15;
				end
				if(in == 4) begin
					state<=4617;
					out<=16;
				end
			end
			2717: begin
				if(in == 0) begin
					state<=2718;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=6607;
					out<=19;
				end
				if(in == 3) begin
					state<=720;
					out<=20;
				end
				if(in == 4) begin
					state<=4618;
					out<=21;
				end
			end
			2718: begin
				if(in == 0) begin
					state<=2719;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=6608;
					out<=24;
				end
				if(in == 3) begin
					state<=721;
					out<=25;
				end
				if(in == 4) begin
					state<=4619;
					out<=26;
				end
			end
			2719: begin
				if(in == 0) begin
					state<=2720;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=6609;
					out<=29;
				end
				if(in == 3) begin
					state<=722;
					out<=30;
				end
				if(in == 4) begin
					state<=4620;
					out<=31;
				end
			end
			2720: begin
				if(in == 0) begin
					state<=2721;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=6610;
					out<=34;
				end
				if(in == 3) begin
					state<=723;
					out<=35;
				end
				if(in == 4) begin
					state<=4621;
					out<=36;
				end
			end
			2721: begin
				if(in == 0) begin
					state<=2722;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=6611;
					out<=39;
				end
				if(in == 3) begin
					state<=724;
					out<=40;
				end
				if(in == 4) begin
					state<=4622;
					out<=41;
				end
			end
			2722: begin
				if(in == 0) begin
					state<=2723;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=6612;
					out<=44;
				end
				if(in == 3) begin
					state<=725;
					out<=45;
				end
				if(in == 4) begin
					state<=4623;
					out<=46;
				end
			end
			2723: begin
				if(in == 0) begin
					state<=2724;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=6613;
					out<=49;
				end
				if(in == 3) begin
					state<=726;
					out<=50;
				end
				if(in == 4) begin
					state<=4624;
					out<=51;
				end
			end
			2724: begin
				if(in == 0) begin
					state<=2725;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=6614;
					out<=54;
				end
				if(in == 3) begin
					state<=727;
					out<=55;
				end
				if(in == 4) begin
					state<=4625;
					out<=56;
				end
			end
			2725: begin
				if(in == 0) begin
					state<=2726;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=6615;
					out<=59;
				end
				if(in == 3) begin
					state<=728;
					out<=60;
				end
				if(in == 4) begin
					state<=4626;
					out<=61;
				end
			end
			2726: begin
				if(in == 0) begin
					state<=2727;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=6616;
					out<=64;
				end
				if(in == 3) begin
					state<=729;
					out<=65;
				end
				if(in == 4) begin
					state<=4627;
					out<=66;
				end
			end
			2727: begin
				if(in == 0) begin
					state<=2728;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=6617;
					out<=69;
				end
				if(in == 3) begin
					state<=730;
					out<=70;
				end
				if(in == 4) begin
					state<=4628;
					out<=71;
				end
			end
			2728: begin
				if(in == 0) begin
					state<=2729;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=6618;
					out<=74;
				end
				if(in == 3) begin
					state<=731;
					out<=75;
				end
				if(in == 4) begin
					state<=4629;
					out<=76;
				end
			end
			2729: begin
				if(in == 0) begin
					state<=2730;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=6619;
					out<=79;
				end
				if(in == 3) begin
					state<=732;
					out<=80;
				end
				if(in == 4) begin
					state<=4630;
					out<=81;
				end
			end
			2730: begin
				if(in == 0) begin
					state<=2731;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=6620;
					out<=84;
				end
				if(in == 3) begin
					state<=733;
					out<=85;
				end
				if(in == 4) begin
					state<=4631;
					out<=86;
				end
			end
			2731: begin
				if(in == 0) begin
					state<=2732;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=6621;
					out<=89;
				end
				if(in == 3) begin
					state<=734;
					out<=90;
				end
				if(in == 4) begin
					state<=4632;
					out<=91;
				end
			end
			2732: begin
				if(in == 0) begin
					state<=2733;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=6622;
					out<=94;
				end
				if(in == 3) begin
					state<=735;
					out<=95;
				end
				if(in == 4) begin
					state<=4633;
					out<=96;
				end
			end
			2733: begin
				if(in == 0) begin
					state<=2734;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=6623;
					out<=99;
				end
				if(in == 3) begin
					state<=736;
					out<=100;
				end
				if(in == 4) begin
					state<=4634;
					out<=101;
				end
			end
			2734: begin
				if(in == 0) begin
					state<=2735;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=6624;
					out<=104;
				end
				if(in == 3) begin
					state<=737;
					out<=105;
				end
				if(in == 4) begin
					state<=4635;
					out<=106;
				end
			end
			2735: begin
				if(in == 0) begin
					state<=2736;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=6625;
					out<=109;
				end
				if(in == 3) begin
					state<=738;
					out<=110;
				end
				if(in == 4) begin
					state<=4636;
					out<=111;
				end
			end
			2736: begin
				if(in == 0) begin
					state<=2737;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=6626;
					out<=114;
				end
				if(in == 3) begin
					state<=739;
					out<=115;
				end
				if(in == 4) begin
					state<=4637;
					out<=116;
				end
			end
			2737: begin
				if(in == 0) begin
					state<=2738;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=6627;
					out<=119;
				end
				if(in == 3) begin
					state<=740;
					out<=120;
				end
				if(in == 4) begin
					state<=4638;
					out<=121;
				end
			end
			2738: begin
				if(in == 0) begin
					state<=2739;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=6628;
					out<=124;
				end
				if(in == 3) begin
					state<=741;
					out<=125;
				end
				if(in == 4) begin
					state<=4639;
					out<=126;
				end
			end
			2739: begin
				if(in == 0) begin
					state<=2740;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=6629;
					out<=129;
				end
				if(in == 3) begin
					state<=742;
					out<=130;
				end
				if(in == 4) begin
					state<=4640;
					out<=131;
				end
			end
			2740: begin
				if(in == 0) begin
					state<=2741;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=6630;
					out<=134;
				end
				if(in == 3) begin
					state<=743;
					out<=135;
				end
				if(in == 4) begin
					state<=4641;
					out<=136;
				end
			end
			2741: begin
				if(in == 0) begin
					state<=2742;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=6631;
					out<=139;
				end
				if(in == 3) begin
					state<=744;
					out<=140;
				end
				if(in == 4) begin
					state<=4642;
					out<=141;
				end
			end
			2742: begin
				if(in == 0) begin
					state<=2743;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=6632;
					out<=144;
				end
				if(in == 3) begin
					state<=745;
					out<=145;
				end
				if(in == 4) begin
					state<=4643;
					out<=146;
				end
			end
			2743: begin
				if(in == 0) begin
					state<=2744;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=6633;
					out<=149;
				end
				if(in == 3) begin
					state<=746;
					out<=150;
				end
				if(in == 4) begin
					state<=4644;
					out<=151;
				end
			end
			2744: begin
				if(in == 0) begin
					state<=2745;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=6634;
					out<=154;
				end
				if(in == 3) begin
					state<=747;
					out<=155;
				end
				if(in == 4) begin
					state<=4645;
					out<=156;
				end
			end
			2745: begin
				if(in == 0) begin
					state<=2746;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=6635;
					out<=159;
				end
				if(in == 3) begin
					state<=748;
					out<=160;
				end
				if(in == 4) begin
					state<=4646;
					out<=161;
				end
			end
			2746: begin
				if(in == 0) begin
					state<=2747;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=6636;
					out<=164;
				end
				if(in == 3) begin
					state<=749;
					out<=165;
				end
				if(in == 4) begin
					state<=4647;
					out<=166;
				end
			end
			2747: begin
				if(in == 0) begin
					state<=2748;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=6637;
					out<=169;
				end
				if(in == 3) begin
					state<=750;
					out<=170;
				end
				if(in == 4) begin
					state<=4648;
					out<=171;
				end
			end
			2748: begin
				if(in == 0) begin
					state<=2749;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=6638;
					out<=174;
				end
				if(in == 3) begin
					state<=751;
					out<=175;
				end
				if(in == 4) begin
					state<=4649;
					out<=176;
				end
			end
			2749: begin
				if(in == 0) begin
					state<=2750;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=6639;
					out<=179;
				end
				if(in == 3) begin
					state<=752;
					out<=180;
				end
				if(in == 4) begin
					state<=4650;
					out<=181;
				end
			end
			2750: begin
				if(in == 0) begin
					state<=2751;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=6640;
					out<=184;
				end
				if(in == 3) begin
					state<=753;
					out<=185;
				end
				if(in == 4) begin
					state<=4651;
					out<=186;
				end
			end
			2751: begin
				if(in == 0) begin
					state<=2752;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=6641;
					out<=189;
				end
				if(in == 3) begin
					state<=754;
					out<=190;
				end
				if(in == 4) begin
					state<=4652;
					out<=191;
				end
			end
			2752: begin
				if(in == 0) begin
					state<=2753;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=6642;
					out<=194;
				end
				if(in == 3) begin
					state<=755;
					out<=195;
				end
				if(in == 4) begin
					state<=4653;
					out<=196;
				end
			end
			2753: begin
				if(in == 0) begin
					state<=2754;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=6643;
					out<=199;
				end
				if(in == 3) begin
					state<=756;
					out<=200;
				end
				if(in == 4) begin
					state<=4654;
					out<=201;
				end
			end
			2754: begin
				if(in == 0) begin
					state<=2755;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=6644;
					out<=204;
				end
				if(in == 3) begin
					state<=757;
					out<=205;
				end
				if(in == 4) begin
					state<=4655;
					out<=206;
				end
			end
			2755: begin
				if(in == 0) begin
					state<=2756;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=6645;
					out<=209;
				end
				if(in == 3) begin
					state<=758;
					out<=210;
				end
				if(in == 4) begin
					state<=4656;
					out<=211;
				end
			end
			2756: begin
				if(in == 0) begin
					state<=2757;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=6646;
					out<=214;
				end
				if(in == 3) begin
					state<=759;
					out<=215;
				end
				if(in == 4) begin
					state<=4657;
					out<=216;
				end
			end
			2757: begin
				if(in == 0) begin
					state<=2758;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=6647;
					out<=219;
				end
				if(in == 3) begin
					state<=760;
					out<=220;
				end
				if(in == 4) begin
					state<=4658;
					out<=221;
				end
			end
			2758: begin
				if(in == 0) begin
					state<=2759;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=6648;
					out<=224;
				end
				if(in == 3) begin
					state<=761;
					out<=225;
				end
				if(in == 4) begin
					state<=4659;
					out<=226;
				end
			end
			2759: begin
				if(in == 0) begin
					state<=2760;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=6649;
					out<=229;
				end
				if(in == 3) begin
					state<=762;
					out<=230;
				end
				if(in == 4) begin
					state<=4660;
					out<=231;
				end
			end
			2760: begin
				if(in == 0) begin
					state<=2761;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=6650;
					out<=234;
				end
				if(in == 3) begin
					state<=763;
					out<=235;
				end
				if(in == 4) begin
					state<=4661;
					out<=236;
				end
			end
			2761: begin
				if(in == 0) begin
					state<=2762;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=6651;
					out<=239;
				end
				if(in == 3) begin
					state<=764;
					out<=240;
				end
				if(in == 4) begin
					state<=4662;
					out<=241;
				end
			end
			2762: begin
				if(in == 0) begin
					state<=2763;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=6652;
					out<=244;
				end
				if(in == 3) begin
					state<=765;
					out<=245;
				end
				if(in == 4) begin
					state<=4663;
					out<=246;
				end
			end
			2763: begin
				if(in == 0) begin
					state<=2764;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=6653;
					out<=249;
				end
				if(in == 3) begin
					state<=766;
					out<=250;
				end
				if(in == 4) begin
					state<=4664;
					out<=251;
				end
			end
			2764: begin
				if(in == 0) begin
					state<=2765;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=6654;
					out<=254;
				end
				if(in == 3) begin
					state<=767;
					out<=255;
				end
				if(in == 4) begin
					state<=4665;
					out<=0;
				end
			end
			2765: begin
				if(in == 0) begin
					state<=2766;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=6655;
					out<=3;
				end
				if(in == 3) begin
					state<=768;
					out<=4;
				end
				if(in == 4) begin
					state<=4666;
					out<=5;
				end
			end
			2766: begin
				if(in == 0) begin
					state<=2767;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=6656;
					out<=8;
				end
				if(in == 3) begin
					state<=769;
					out<=9;
				end
				if(in == 4) begin
					state<=4667;
					out<=10;
				end
			end
			2767: begin
				if(in == 0) begin
					state<=2768;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=6657;
					out<=13;
				end
				if(in == 3) begin
					state<=770;
					out<=14;
				end
				if(in == 4) begin
					state<=4668;
					out<=15;
				end
			end
			2768: begin
				if(in == 0) begin
					state<=2769;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=6658;
					out<=18;
				end
				if(in == 3) begin
					state<=771;
					out<=19;
				end
				if(in == 4) begin
					state<=4669;
					out<=20;
				end
			end
			2769: begin
				if(in == 0) begin
					state<=2770;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=6659;
					out<=23;
				end
				if(in == 3) begin
					state<=772;
					out<=24;
				end
				if(in == 4) begin
					state<=4670;
					out<=25;
				end
			end
			2770: begin
				if(in == 0) begin
					state<=2771;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=6660;
					out<=28;
				end
				if(in == 3) begin
					state<=773;
					out<=29;
				end
				if(in == 4) begin
					state<=4671;
					out<=30;
				end
			end
			2771: begin
				if(in == 0) begin
					state<=2772;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=6661;
					out<=33;
				end
				if(in == 3) begin
					state<=774;
					out<=34;
				end
				if(in == 4) begin
					state<=4672;
					out<=35;
				end
			end
			2772: begin
				if(in == 0) begin
					state<=2773;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=6662;
					out<=38;
				end
				if(in == 3) begin
					state<=775;
					out<=39;
				end
				if(in == 4) begin
					state<=4673;
					out<=40;
				end
			end
			2773: begin
				if(in == 0) begin
					state<=2774;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=6663;
					out<=43;
				end
				if(in == 3) begin
					state<=776;
					out<=44;
				end
				if(in == 4) begin
					state<=4674;
					out<=45;
				end
			end
			2774: begin
				if(in == 0) begin
					state<=2775;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=6664;
					out<=48;
				end
				if(in == 3) begin
					state<=777;
					out<=49;
				end
				if(in == 4) begin
					state<=4675;
					out<=50;
				end
			end
			2775: begin
				if(in == 0) begin
					state<=2776;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=6665;
					out<=53;
				end
				if(in == 3) begin
					state<=778;
					out<=54;
				end
				if(in == 4) begin
					state<=4676;
					out<=55;
				end
			end
			2776: begin
				if(in == 0) begin
					state<=2777;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=6666;
					out<=58;
				end
				if(in == 3) begin
					state<=779;
					out<=59;
				end
				if(in == 4) begin
					state<=4677;
					out<=60;
				end
			end
			2777: begin
				if(in == 0) begin
					state<=2778;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=6667;
					out<=63;
				end
				if(in == 3) begin
					state<=780;
					out<=64;
				end
				if(in == 4) begin
					state<=4678;
					out<=65;
				end
			end
			2778: begin
				if(in == 0) begin
					state<=2779;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=6668;
					out<=68;
				end
				if(in == 3) begin
					state<=781;
					out<=69;
				end
				if(in == 4) begin
					state<=4679;
					out<=70;
				end
			end
			2779: begin
				if(in == 0) begin
					state<=2780;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=6669;
					out<=73;
				end
				if(in == 3) begin
					state<=782;
					out<=74;
				end
				if(in == 4) begin
					state<=4680;
					out<=75;
				end
			end
			2780: begin
				if(in == 0) begin
					state<=2781;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=6670;
					out<=78;
				end
				if(in == 3) begin
					state<=783;
					out<=79;
				end
				if(in == 4) begin
					state<=4681;
					out<=80;
				end
			end
			2781: begin
				if(in == 0) begin
					state<=2782;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=6671;
					out<=83;
				end
				if(in == 3) begin
					state<=784;
					out<=84;
				end
				if(in == 4) begin
					state<=4682;
					out<=85;
				end
			end
			2782: begin
				if(in == 0) begin
					state<=2783;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=6672;
					out<=88;
				end
				if(in == 3) begin
					state<=785;
					out<=89;
				end
				if(in == 4) begin
					state<=4683;
					out<=90;
				end
			end
			2783: begin
				if(in == 0) begin
					state<=2784;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=6673;
					out<=93;
				end
				if(in == 3) begin
					state<=786;
					out<=94;
				end
				if(in == 4) begin
					state<=4684;
					out<=95;
				end
			end
			2784: begin
				if(in == 0) begin
					state<=2785;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=6674;
					out<=98;
				end
				if(in == 3) begin
					state<=787;
					out<=99;
				end
				if(in == 4) begin
					state<=4685;
					out<=100;
				end
			end
			2785: begin
				if(in == 0) begin
					state<=2786;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=6675;
					out<=103;
				end
				if(in == 3) begin
					state<=788;
					out<=104;
				end
				if(in == 4) begin
					state<=4686;
					out<=105;
				end
			end
			2786: begin
				if(in == 0) begin
					state<=2787;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=6676;
					out<=108;
				end
				if(in == 3) begin
					state<=789;
					out<=109;
				end
				if(in == 4) begin
					state<=4687;
					out<=110;
				end
			end
			2787: begin
				if(in == 0) begin
					state<=2788;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=6677;
					out<=113;
				end
				if(in == 3) begin
					state<=790;
					out<=114;
				end
				if(in == 4) begin
					state<=4688;
					out<=115;
				end
			end
			2788: begin
				if(in == 0) begin
					state<=2789;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=6678;
					out<=118;
				end
				if(in == 3) begin
					state<=791;
					out<=119;
				end
				if(in == 4) begin
					state<=4689;
					out<=120;
				end
			end
			2789: begin
				if(in == 0) begin
					state<=2790;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=6679;
					out<=123;
				end
				if(in == 3) begin
					state<=792;
					out<=124;
				end
				if(in == 4) begin
					state<=4690;
					out<=125;
				end
			end
			2790: begin
				if(in == 0) begin
					state<=2791;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=6680;
					out<=128;
				end
				if(in == 3) begin
					state<=793;
					out<=129;
				end
				if(in == 4) begin
					state<=4691;
					out<=130;
				end
			end
			2791: begin
				if(in == 0) begin
					state<=2792;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=6681;
					out<=133;
				end
				if(in == 3) begin
					state<=794;
					out<=134;
				end
				if(in == 4) begin
					state<=4692;
					out<=135;
				end
			end
			2792: begin
				if(in == 0) begin
					state<=2793;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=6682;
					out<=138;
				end
				if(in == 3) begin
					state<=795;
					out<=139;
				end
				if(in == 4) begin
					state<=4693;
					out<=140;
				end
			end
			2793: begin
				if(in == 0) begin
					state<=2794;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=6683;
					out<=143;
				end
				if(in == 3) begin
					state<=796;
					out<=144;
				end
				if(in == 4) begin
					state<=4694;
					out<=145;
				end
			end
			2794: begin
				if(in == 0) begin
					state<=2795;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=6684;
					out<=148;
				end
				if(in == 3) begin
					state<=797;
					out<=149;
				end
				if(in == 4) begin
					state<=4695;
					out<=150;
				end
			end
			2795: begin
				if(in == 0) begin
					state<=2796;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=6685;
					out<=153;
				end
				if(in == 3) begin
					state<=798;
					out<=154;
				end
				if(in == 4) begin
					state<=4696;
					out<=155;
				end
			end
			2796: begin
				if(in == 0) begin
					state<=2797;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=6686;
					out<=158;
				end
				if(in == 3) begin
					state<=799;
					out<=159;
				end
				if(in == 4) begin
					state<=4697;
					out<=160;
				end
			end
			2797: begin
				if(in == 0) begin
					state<=2808;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=6697;
					out<=163;
				end
				if(in == 3) begin
					state<=810;
					out<=164;
				end
				if(in == 4) begin
					state<=4708;
					out<=165;
				end
			end
			2798: begin
				if(in == 0) begin
					state<=2799;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=6688;
					out<=168;
				end
				if(in == 3) begin
					state<=801;
					out<=169;
				end
				if(in == 4) begin
					state<=4699;
					out<=170;
				end
			end
			2799: begin
				if(in == 0) begin
					state<=2800;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=6689;
					out<=173;
				end
				if(in == 3) begin
					state<=802;
					out<=174;
				end
				if(in == 4) begin
					state<=4700;
					out<=175;
				end
			end
			2800: begin
				if(in == 0) begin
					state<=2801;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=6690;
					out<=178;
				end
				if(in == 3) begin
					state<=803;
					out<=179;
				end
				if(in == 4) begin
					state<=4701;
					out<=180;
				end
			end
			2801: begin
				if(in == 0) begin
					state<=2802;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=6691;
					out<=183;
				end
				if(in == 3) begin
					state<=804;
					out<=184;
				end
				if(in == 4) begin
					state<=4702;
					out<=185;
				end
			end
			2802: begin
				if(in == 0) begin
					state<=2803;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=6692;
					out<=188;
				end
				if(in == 3) begin
					state<=805;
					out<=189;
				end
				if(in == 4) begin
					state<=4703;
					out<=190;
				end
			end
			2803: begin
				if(in == 0) begin
					state<=2804;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=6693;
					out<=193;
				end
				if(in == 3) begin
					state<=806;
					out<=194;
				end
				if(in == 4) begin
					state<=4704;
					out<=195;
				end
			end
			2804: begin
				if(in == 0) begin
					state<=2805;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=6694;
					out<=198;
				end
				if(in == 3) begin
					state<=807;
					out<=199;
				end
				if(in == 4) begin
					state<=4705;
					out<=200;
				end
			end
			2805: begin
				if(in == 0) begin
					state<=2806;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=6695;
					out<=203;
				end
				if(in == 3) begin
					state<=808;
					out<=204;
				end
				if(in == 4) begin
					state<=4706;
					out<=205;
				end
			end
			2806: begin
				if(in == 0) begin
					state<=2807;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=6696;
					out<=208;
				end
				if(in == 3) begin
					state<=809;
					out<=209;
				end
				if(in == 4) begin
					state<=4707;
					out<=210;
				end
			end
			2807: begin
				if(in == 0) begin
					state<=3509;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=7398;
					out<=213;
				end
				if(in == 3) begin
					state<=1608;
					out<=214;
				end
				if(in == 4) begin
					state<=5497;
					out<=215;
				end
			end
			2808: begin
				if(in == 0) begin
					state<=2809;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=6698;
					out<=218;
				end
				if(in == 3) begin
					state<=811;
					out<=219;
				end
				if(in == 4) begin
					state<=4709;
					out<=220;
				end
			end
			2809: begin
				if(in == 0) begin
					state<=2810;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=6699;
					out<=223;
				end
				if(in == 3) begin
					state<=812;
					out<=224;
				end
				if(in == 4) begin
					state<=4710;
					out<=225;
				end
			end
			2810: begin
				if(in == 0) begin
					state<=2811;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=6700;
					out<=228;
				end
				if(in == 3) begin
					state<=813;
					out<=229;
				end
				if(in == 4) begin
					state<=4711;
					out<=230;
				end
			end
			2811: begin
				if(in == 0) begin
					state<=2812;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=6701;
					out<=233;
				end
				if(in == 3) begin
					state<=814;
					out<=234;
				end
				if(in == 4) begin
					state<=4712;
					out<=235;
				end
			end
			2812: begin
				if(in == 0) begin
					state<=2813;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=6702;
					out<=238;
				end
				if(in == 3) begin
					state<=815;
					out<=239;
				end
				if(in == 4) begin
					state<=4713;
					out<=240;
				end
			end
			2813: begin
				if(in == 0) begin
					state<=2814;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=6703;
					out<=243;
				end
				if(in == 3) begin
					state<=816;
					out<=244;
				end
				if(in == 4) begin
					state<=4714;
					out<=245;
				end
			end
			2814: begin
				if(in == 0) begin
					state<=2815;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=6704;
					out<=248;
				end
				if(in == 3) begin
					state<=817;
					out<=249;
				end
				if(in == 4) begin
					state<=4715;
					out<=250;
				end
			end
			2815: begin
				if(in == 0) begin
					state<=2816;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=6705;
					out<=253;
				end
				if(in == 3) begin
					state<=818;
					out<=254;
				end
				if(in == 4) begin
					state<=4716;
					out<=255;
				end
			end
			2816: begin
				if(in == 0) begin
					state<=2817;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=6706;
					out<=2;
				end
				if(in == 3) begin
					state<=819;
					out<=3;
				end
				if(in == 4) begin
					state<=4717;
					out<=4;
				end
			end
			2817: begin
				if(in == 0) begin
					state<=2818;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=6707;
					out<=7;
				end
				if(in == 3) begin
					state<=820;
					out<=8;
				end
				if(in == 4) begin
					state<=4718;
					out<=9;
				end
			end
			2818: begin
				if(in == 0) begin
					state<=2819;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=6708;
					out<=12;
				end
				if(in == 3) begin
					state<=821;
					out<=13;
				end
				if(in == 4) begin
					state<=4719;
					out<=14;
				end
			end
			2819: begin
				if(in == 0) begin
					state<=2820;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=6709;
					out<=17;
				end
				if(in == 3) begin
					state<=822;
					out<=18;
				end
				if(in == 4) begin
					state<=4720;
					out<=19;
				end
			end
			2820: begin
				if(in == 0) begin
					state<=2821;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=6710;
					out<=22;
				end
				if(in == 3) begin
					state<=823;
					out<=23;
				end
				if(in == 4) begin
					state<=4721;
					out<=24;
				end
			end
			2821: begin
				if(in == 0) begin
					state<=2822;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=6711;
					out<=27;
				end
				if(in == 3) begin
					state<=824;
					out<=28;
				end
				if(in == 4) begin
					state<=4722;
					out<=29;
				end
			end
			2822: begin
				if(in == 0) begin
					state<=2823;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=6712;
					out<=32;
				end
				if(in == 3) begin
					state<=825;
					out<=33;
				end
				if(in == 4) begin
					state<=4723;
					out<=34;
				end
			end
			2823: begin
				if(in == 0) begin
					state<=2824;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=6713;
					out<=37;
				end
				if(in == 3) begin
					state<=826;
					out<=38;
				end
				if(in == 4) begin
					state<=4724;
					out<=39;
				end
			end
			2824: begin
				if(in == 0) begin
					state<=2825;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=6714;
					out<=42;
				end
				if(in == 3) begin
					state<=827;
					out<=43;
				end
				if(in == 4) begin
					state<=4725;
					out<=44;
				end
			end
			2825: begin
				if(in == 0) begin
					state<=2826;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=6715;
					out<=47;
				end
				if(in == 3) begin
					state<=828;
					out<=48;
				end
				if(in == 4) begin
					state<=4726;
					out<=49;
				end
			end
			2826: begin
				if(in == 0) begin
					state<=2827;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=6716;
					out<=52;
				end
				if(in == 3) begin
					state<=829;
					out<=53;
				end
				if(in == 4) begin
					state<=4727;
					out<=54;
				end
			end
			2827: begin
				if(in == 0) begin
					state<=2828;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=6717;
					out<=57;
				end
				if(in == 3) begin
					state<=830;
					out<=58;
				end
				if(in == 4) begin
					state<=4728;
					out<=59;
				end
			end
			2828: begin
				if(in == 0) begin
					state<=2829;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=6718;
					out<=62;
				end
				if(in == 3) begin
					state<=831;
					out<=63;
				end
				if(in == 4) begin
					state<=4729;
					out<=64;
				end
			end
			2829: begin
				if(in == 0) begin
					state<=2830;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=6719;
					out<=67;
				end
				if(in == 3) begin
					state<=832;
					out<=68;
				end
				if(in == 4) begin
					state<=4730;
					out<=69;
				end
			end
			2830: begin
				if(in == 0) begin
					state<=2831;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=6720;
					out<=72;
				end
				if(in == 3) begin
					state<=833;
					out<=73;
				end
				if(in == 4) begin
					state<=4731;
					out<=74;
				end
			end
			2831: begin
				if(in == 0) begin
					state<=2832;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=6721;
					out<=77;
				end
				if(in == 3) begin
					state<=834;
					out<=78;
				end
				if(in == 4) begin
					state<=4732;
					out<=79;
				end
			end
			2832: begin
				if(in == 0) begin
					state<=2833;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=6722;
					out<=82;
				end
				if(in == 3) begin
					state<=835;
					out<=83;
				end
				if(in == 4) begin
					state<=4733;
					out<=84;
				end
			end
			2833: begin
				if(in == 0) begin
					state<=2834;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=6723;
					out<=87;
				end
				if(in == 3) begin
					state<=836;
					out<=88;
				end
				if(in == 4) begin
					state<=4734;
					out<=89;
				end
			end
			2834: begin
				if(in == 0) begin
					state<=2835;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=6724;
					out<=92;
				end
				if(in == 3) begin
					state<=837;
					out<=93;
				end
				if(in == 4) begin
					state<=4735;
					out<=94;
				end
			end
			2835: begin
				if(in == 0) begin
					state<=2836;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=6725;
					out<=97;
				end
				if(in == 3) begin
					state<=838;
					out<=98;
				end
				if(in == 4) begin
					state<=4736;
					out<=99;
				end
			end
			2836: begin
				if(in == 0) begin
					state<=2837;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=6726;
					out<=102;
				end
				if(in == 3) begin
					state<=839;
					out<=103;
				end
				if(in == 4) begin
					state<=4737;
					out<=104;
				end
			end
			2837: begin
				if(in == 0) begin
					state<=2838;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=6727;
					out<=107;
				end
				if(in == 3) begin
					state<=840;
					out<=108;
				end
				if(in == 4) begin
					state<=4738;
					out<=109;
				end
			end
			2838: begin
				if(in == 0) begin
					state<=2839;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=6728;
					out<=112;
				end
				if(in == 3) begin
					state<=841;
					out<=113;
				end
				if(in == 4) begin
					state<=4739;
					out<=114;
				end
			end
			2839: begin
				if(in == 0) begin
					state<=2840;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=6729;
					out<=117;
				end
				if(in == 3) begin
					state<=842;
					out<=118;
				end
				if(in == 4) begin
					state<=4740;
					out<=119;
				end
			end
			2840: begin
				if(in == 0) begin
					state<=2841;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=6730;
					out<=122;
				end
				if(in == 3) begin
					state<=843;
					out<=123;
				end
				if(in == 4) begin
					state<=4741;
					out<=124;
				end
			end
			2841: begin
				if(in == 0) begin
					state<=2842;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=6731;
					out<=127;
				end
				if(in == 3) begin
					state<=844;
					out<=128;
				end
				if(in == 4) begin
					state<=4742;
					out<=129;
				end
			end
			2842: begin
				if(in == 0) begin
					state<=2843;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=6732;
					out<=132;
				end
				if(in == 3) begin
					state<=845;
					out<=133;
				end
				if(in == 4) begin
					state<=4743;
					out<=134;
				end
			end
			2843: begin
				if(in == 0) begin
					state<=2844;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=6733;
					out<=137;
				end
				if(in == 3) begin
					state<=846;
					out<=138;
				end
				if(in == 4) begin
					state<=4744;
					out<=139;
				end
			end
			2844: begin
				if(in == 0) begin
					state<=2845;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=6734;
					out<=142;
				end
				if(in == 3) begin
					state<=847;
					out<=143;
				end
				if(in == 4) begin
					state<=4745;
					out<=144;
				end
			end
			2845: begin
				if(in == 0) begin
					state<=2846;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=6735;
					out<=147;
				end
				if(in == 3) begin
					state<=848;
					out<=148;
				end
				if(in == 4) begin
					state<=4746;
					out<=149;
				end
			end
			2846: begin
				if(in == 0) begin
					state<=2847;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=6736;
					out<=152;
				end
				if(in == 3) begin
					state<=849;
					out<=153;
				end
				if(in == 4) begin
					state<=4747;
					out<=154;
				end
			end
			2847: begin
				if(in == 0) begin
					state<=2848;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=6737;
					out<=157;
				end
				if(in == 3) begin
					state<=850;
					out<=158;
				end
				if(in == 4) begin
					state<=4748;
					out<=159;
				end
			end
			2848: begin
				if(in == 0) begin
					state<=2849;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=6738;
					out<=162;
				end
				if(in == 3) begin
					state<=851;
					out<=163;
				end
				if(in == 4) begin
					state<=4749;
					out<=164;
				end
			end
			2849: begin
				if(in == 0) begin
					state<=2850;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=6739;
					out<=167;
				end
				if(in == 3) begin
					state<=852;
					out<=168;
				end
				if(in == 4) begin
					state<=4750;
					out<=169;
				end
			end
			2850: begin
				if(in == 0) begin
					state<=2851;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=6740;
					out<=172;
				end
				if(in == 3) begin
					state<=853;
					out<=173;
				end
				if(in == 4) begin
					state<=4751;
					out<=174;
				end
			end
			2851: begin
				if(in == 0) begin
					state<=2852;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=6741;
					out<=177;
				end
				if(in == 3) begin
					state<=854;
					out<=178;
				end
				if(in == 4) begin
					state<=4752;
					out<=179;
				end
			end
			2852: begin
				if(in == 0) begin
					state<=2853;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=6742;
					out<=182;
				end
				if(in == 3) begin
					state<=855;
					out<=183;
				end
				if(in == 4) begin
					state<=4753;
					out<=184;
				end
			end
			2853: begin
				if(in == 0) begin
					state<=2854;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=6743;
					out<=187;
				end
				if(in == 3) begin
					state<=856;
					out<=188;
				end
				if(in == 4) begin
					state<=4754;
					out<=189;
				end
			end
			2854: begin
				if(in == 0) begin
					state<=2855;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=6744;
					out<=192;
				end
				if(in == 3) begin
					state<=857;
					out<=193;
				end
				if(in == 4) begin
					state<=4755;
					out<=194;
				end
			end
			2855: begin
				if(in == 0) begin
					state<=2856;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=6745;
					out<=197;
				end
				if(in == 3) begin
					state<=858;
					out<=198;
				end
				if(in == 4) begin
					state<=4756;
					out<=199;
				end
			end
			2856: begin
				if(in == 0) begin
					state<=2857;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=6746;
					out<=202;
				end
				if(in == 3) begin
					state<=859;
					out<=203;
				end
				if(in == 4) begin
					state<=4757;
					out<=204;
				end
			end
			2857: begin
				if(in == 0) begin
					state<=2858;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=6747;
					out<=207;
				end
				if(in == 3) begin
					state<=860;
					out<=208;
				end
				if(in == 4) begin
					state<=4758;
					out<=209;
				end
			end
			2858: begin
				if(in == 0) begin
					state<=2859;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=6748;
					out<=212;
				end
				if(in == 3) begin
					state<=861;
					out<=213;
				end
				if(in == 4) begin
					state<=4759;
					out<=214;
				end
			end
			2859: begin
				if(in == 0) begin
					state<=2860;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=6749;
					out<=217;
				end
				if(in == 3) begin
					state<=862;
					out<=218;
				end
				if(in == 4) begin
					state<=4760;
					out<=219;
				end
			end
			2860: begin
				if(in == 0) begin
					state<=2861;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=6750;
					out<=222;
				end
				if(in == 3) begin
					state<=863;
					out<=223;
				end
				if(in == 4) begin
					state<=4761;
					out<=224;
				end
			end
			2861: begin
				if(in == 0) begin
					state<=2862;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=6751;
					out<=227;
				end
				if(in == 3) begin
					state<=864;
					out<=228;
				end
				if(in == 4) begin
					state<=4762;
					out<=229;
				end
			end
			2862: begin
				if(in == 0) begin
					state<=2863;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=6752;
					out<=232;
				end
				if(in == 3) begin
					state<=865;
					out<=233;
				end
				if(in == 4) begin
					state<=4763;
					out<=234;
				end
			end
			2863: begin
				if(in == 0) begin
					state<=2864;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=6753;
					out<=237;
				end
				if(in == 3) begin
					state<=866;
					out<=238;
				end
				if(in == 4) begin
					state<=4764;
					out<=239;
				end
			end
			2864: begin
				if(in == 0) begin
					state<=2865;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=6754;
					out<=242;
				end
				if(in == 3) begin
					state<=867;
					out<=243;
				end
				if(in == 4) begin
					state<=4765;
					out<=244;
				end
			end
			2865: begin
				if(in == 0) begin
					state<=2866;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=6755;
					out<=247;
				end
				if(in == 3) begin
					state<=868;
					out<=248;
				end
				if(in == 4) begin
					state<=4766;
					out<=249;
				end
			end
			2866: begin
				if(in == 0) begin
					state<=2867;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=6756;
					out<=252;
				end
				if(in == 3) begin
					state<=869;
					out<=253;
				end
				if(in == 4) begin
					state<=4767;
					out<=254;
				end
			end
			2867: begin
				if(in == 0) begin
					state<=2868;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=6757;
					out<=1;
				end
				if(in == 3) begin
					state<=870;
					out<=2;
				end
				if(in == 4) begin
					state<=4768;
					out<=3;
				end
			end
			2868: begin
				if(in == 0) begin
					state<=2869;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=6758;
					out<=6;
				end
				if(in == 3) begin
					state<=871;
					out<=7;
				end
				if(in == 4) begin
					state<=4769;
					out<=8;
				end
			end
			2869: begin
				if(in == 0) begin
					state<=2870;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=6759;
					out<=11;
				end
				if(in == 3) begin
					state<=872;
					out<=12;
				end
				if(in == 4) begin
					state<=4770;
					out<=13;
				end
			end
			2870: begin
				if(in == 0) begin
					state<=2871;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=6760;
					out<=16;
				end
				if(in == 3) begin
					state<=873;
					out<=17;
				end
				if(in == 4) begin
					state<=4771;
					out<=18;
				end
			end
			2871: begin
				if(in == 0) begin
					state<=2872;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=6761;
					out<=21;
				end
				if(in == 3) begin
					state<=874;
					out<=22;
				end
				if(in == 4) begin
					state<=4772;
					out<=23;
				end
			end
			2872: begin
				if(in == 0) begin
					state<=2873;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=6762;
					out<=26;
				end
				if(in == 3) begin
					state<=875;
					out<=27;
				end
				if(in == 4) begin
					state<=4773;
					out<=28;
				end
			end
			2873: begin
				if(in == 0) begin
					state<=2874;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=6763;
					out<=31;
				end
				if(in == 3) begin
					state<=876;
					out<=32;
				end
				if(in == 4) begin
					state<=4774;
					out<=33;
				end
			end
			2874: begin
				if(in == 0) begin
					state<=2875;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=6764;
					out<=36;
				end
				if(in == 3) begin
					state<=877;
					out<=37;
				end
				if(in == 4) begin
					state<=4775;
					out<=38;
				end
			end
			2875: begin
				if(in == 0) begin
					state<=2876;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=6765;
					out<=41;
				end
				if(in == 3) begin
					state<=878;
					out<=42;
				end
				if(in == 4) begin
					state<=4776;
					out<=43;
				end
			end
			2876: begin
				if(in == 0) begin
					state<=2877;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=6766;
					out<=46;
				end
				if(in == 3) begin
					state<=879;
					out<=47;
				end
				if(in == 4) begin
					state<=4777;
					out<=48;
				end
			end
			2877: begin
				if(in == 0) begin
					state<=2878;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=6767;
					out<=51;
				end
				if(in == 3) begin
					state<=880;
					out<=52;
				end
				if(in == 4) begin
					state<=4778;
					out<=53;
				end
			end
			2878: begin
				if(in == 0) begin
					state<=2879;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=6768;
					out<=56;
				end
				if(in == 3) begin
					state<=881;
					out<=57;
				end
				if(in == 4) begin
					state<=4779;
					out<=58;
				end
			end
			2879: begin
				if(in == 0) begin
					state<=2880;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=6769;
					out<=61;
				end
				if(in == 3) begin
					state<=882;
					out<=62;
				end
				if(in == 4) begin
					state<=4780;
					out<=63;
				end
			end
			2880: begin
				if(in == 0) begin
					state<=2881;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=6770;
					out<=66;
				end
				if(in == 3) begin
					state<=883;
					out<=67;
				end
				if(in == 4) begin
					state<=4781;
					out<=68;
				end
			end
			2881: begin
				if(in == 0) begin
					state<=2882;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=6771;
					out<=71;
				end
				if(in == 3) begin
					state<=884;
					out<=72;
				end
				if(in == 4) begin
					state<=4782;
					out<=73;
				end
			end
			2882: begin
				if(in == 0) begin
					state<=2883;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=6772;
					out<=76;
				end
				if(in == 3) begin
					state<=885;
					out<=77;
				end
				if(in == 4) begin
					state<=4783;
					out<=78;
				end
			end
			2883: begin
				if(in == 0) begin
					state<=2884;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=6773;
					out<=81;
				end
				if(in == 3) begin
					state<=886;
					out<=82;
				end
				if(in == 4) begin
					state<=4784;
					out<=83;
				end
			end
			2884: begin
				if(in == 0) begin
					state<=2885;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=6774;
					out<=86;
				end
				if(in == 3) begin
					state<=887;
					out<=87;
				end
				if(in == 4) begin
					state<=4785;
					out<=88;
				end
			end
			2885: begin
				if(in == 0) begin
					state<=2886;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=6775;
					out<=91;
				end
				if(in == 3) begin
					state<=888;
					out<=92;
				end
				if(in == 4) begin
					state<=4786;
					out<=93;
				end
			end
			2886: begin
				if(in == 0) begin
					state<=2887;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=6776;
					out<=96;
				end
				if(in == 3) begin
					state<=889;
					out<=97;
				end
				if(in == 4) begin
					state<=4787;
					out<=98;
				end
			end
			2887: begin
				if(in == 0) begin
					state<=2888;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=6777;
					out<=101;
				end
				if(in == 3) begin
					state<=890;
					out<=102;
				end
				if(in == 4) begin
					state<=4788;
					out<=103;
				end
			end
			2888: begin
				if(in == 0) begin
					state<=2889;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=6778;
					out<=106;
				end
				if(in == 3) begin
					state<=891;
					out<=107;
				end
				if(in == 4) begin
					state<=4789;
					out<=108;
				end
			end
			2889: begin
				if(in == 0) begin
					state<=2890;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=6779;
					out<=111;
				end
				if(in == 3) begin
					state<=892;
					out<=112;
				end
				if(in == 4) begin
					state<=4790;
					out<=113;
				end
			end
			2890: begin
				if(in == 0) begin
					state<=2891;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=6780;
					out<=116;
				end
				if(in == 3) begin
					state<=893;
					out<=117;
				end
				if(in == 4) begin
					state<=4791;
					out<=118;
				end
			end
			2891: begin
				if(in == 0) begin
					state<=2892;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=6781;
					out<=121;
				end
				if(in == 3) begin
					state<=894;
					out<=122;
				end
				if(in == 4) begin
					state<=4792;
					out<=123;
				end
			end
			2892: begin
				if(in == 0) begin
					state<=2893;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=6782;
					out<=126;
				end
				if(in == 3) begin
					state<=895;
					out<=127;
				end
				if(in == 4) begin
					state<=4793;
					out<=128;
				end
			end
			2893: begin
				if(in == 0) begin
					state<=2894;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=6783;
					out<=131;
				end
				if(in == 3) begin
					state<=896;
					out<=132;
				end
				if(in == 4) begin
					state<=4794;
					out<=133;
				end
			end
			2894: begin
				if(in == 0) begin
					state<=2895;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=6784;
					out<=136;
				end
				if(in == 3) begin
					state<=897;
					out<=137;
				end
				if(in == 4) begin
					state<=4795;
					out<=138;
				end
			end
			2895: begin
				if(in == 0) begin
					state<=2896;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=6785;
					out<=141;
				end
				if(in == 3) begin
					state<=898;
					out<=142;
				end
				if(in == 4) begin
					state<=4796;
					out<=143;
				end
			end
			2896: begin
				if(in == 0) begin
					state<=2897;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=6786;
					out<=146;
				end
				if(in == 3) begin
					state<=899;
					out<=147;
				end
				if(in == 4) begin
					state<=4797;
					out<=148;
				end
			end
			2897: begin
				if(in == 0) begin
					state<=2798;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=6687;
					out<=151;
				end
				if(in == 3) begin
					state<=800;
					out<=152;
				end
				if(in == 4) begin
					state<=4698;
					out<=153;
				end
			end
			2898: begin
				if(in == 0) begin
					state<=2899;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=6788;
					out<=156;
				end
				if(in == 3) begin
					state<=1454;
					out<=157;
				end
				if(in == 4) begin
					state<=5343;
					out<=158;
				end
			end
			2899: begin
				if(in == 0) begin
					state<=2900;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=6789;
					out<=161;
				end
				if(in == 3) begin
					state<=1455;
					out<=162;
				end
				if(in == 4) begin
					state<=5344;
					out<=163;
				end
			end
			2900: begin
				if(in == 0) begin
					state<=2901;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=6790;
					out<=166;
				end
				if(in == 3) begin
					state<=1456;
					out<=167;
				end
				if(in == 4) begin
					state<=5345;
					out<=168;
				end
			end
			2901: begin
				if(in == 0) begin
					state<=2902;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=6791;
					out<=171;
				end
				if(in == 3) begin
					state<=1457;
					out<=172;
				end
				if(in == 4) begin
					state<=5346;
					out<=173;
				end
			end
			2902: begin
				if(in == 0) begin
					state<=2903;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=6792;
					out<=176;
				end
				if(in == 3) begin
					state<=1458;
					out<=177;
				end
				if(in == 4) begin
					state<=5347;
					out<=178;
				end
			end
			2903: begin
				if(in == 0) begin
					state<=2904;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=6793;
					out<=181;
				end
				if(in == 3) begin
					state<=1459;
					out<=182;
				end
				if(in == 4) begin
					state<=5348;
					out<=183;
				end
			end
			2904: begin
				if(in == 0) begin
					state<=2905;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=6794;
					out<=186;
				end
				if(in == 3) begin
					state<=1460;
					out<=187;
				end
				if(in == 4) begin
					state<=5349;
					out<=188;
				end
			end
			2905: begin
				if(in == 0) begin
					state<=2906;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=6795;
					out<=191;
				end
				if(in == 3) begin
					state<=1461;
					out<=192;
				end
				if(in == 4) begin
					state<=5350;
					out<=193;
				end
			end
			2906: begin
				if(in == 0) begin
					state<=2907;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=6796;
					out<=196;
				end
				if(in == 3) begin
					state<=1462;
					out<=197;
				end
				if(in == 4) begin
					state<=5351;
					out<=198;
				end
			end
			2907: begin
				if(in == 0) begin
					state<=2908;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=6797;
					out<=201;
				end
				if(in == 3) begin
					state<=1463;
					out<=202;
				end
				if(in == 4) begin
					state<=5352;
					out<=203;
				end
			end
			2908: begin
				if(in == 0) begin
					state<=2909;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=6798;
					out<=206;
				end
				if(in == 3) begin
					state<=1464;
					out<=207;
				end
				if(in == 4) begin
					state<=5353;
					out<=208;
				end
			end
			2909: begin
				if(in == 0) begin
					state<=2910;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=6799;
					out<=211;
				end
				if(in == 3) begin
					state<=1465;
					out<=212;
				end
				if(in == 4) begin
					state<=5354;
					out<=213;
				end
			end
			2910: begin
				if(in == 0) begin
					state<=2911;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=6800;
					out<=216;
				end
				if(in == 3) begin
					state<=1466;
					out<=217;
				end
				if(in == 4) begin
					state<=5355;
					out<=218;
				end
			end
			2911: begin
				if(in == 0) begin
					state<=2912;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=6801;
					out<=221;
				end
				if(in == 3) begin
					state<=1467;
					out<=222;
				end
				if(in == 4) begin
					state<=5356;
					out<=223;
				end
			end
			2912: begin
				if(in == 0) begin
					state<=2913;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=6802;
					out<=226;
				end
				if(in == 3) begin
					state<=1468;
					out<=227;
				end
				if(in == 4) begin
					state<=5357;
					out<=228;
				end
			end
			2913: begin
				if(in == 0) begin
					state<=2914;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=6803;
					out<=231;
				end
				if(in == 3) begin
					state<=1469;
					out<=232;
				end
				if(in == 4) begin
					state<=5358;
					out<=233;
				end
			end
			2914: begin
				if(in == 0) begin
					state<=2915;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=6804;
					out<=236;
				end
				if(in == 3) begin
					state<=1470;
					out<=237;
				end
				if(in == 4) begin
					state<=5359;
					out<=238;
				end
			end
			2915: begin
				if(in == 0) begin
					state<=2916;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=6805;
					out<=241;
				end
				if(in == 3) begin
					state<=1471;
					out<=242;
				end
				if(in == 4) begin
					state<=5360;
					out<=243;
				end
			end
			2916: begin
				if(in == 0) begin
					state<=2917;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=6806;
					out<=246;
				end
				if(in == 3) begin
					state<=1472;
					out<=247;
				end
				if(in == 4) begin
					state<=5361;
					out<=248;
				end
			end
			2917: begin
				if(in == 0) begin
					state<=2918;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=6807;
					out<=251;
				end
				if(in == 3) begin
					state<=1473;
					out<=252;
				end
				if(in == 4) begin
					state<=5362;
					out<=253;
				end
			end
			2918: begin
				if(in == 0) begin
					state<=2919;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=6808;
					out<=0;
				end
				if(in == 3) begin
					state<=1474;
					out<=1;
				end
				if(in == 4) begin
					state<=5363;
					out<=2;
				end
			end
			2919: begin
				if(in == 0) begin
					state<=2920;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=6809;
					out<=5;
				end
				if(in == 3) begin
					state<=1475;
					out<=6;
				end
				if(in == 4) begin
					state<=5364;
					out<=7;
				end
			end
			2920: begin
				if(in == 0) begin
					state<=2921;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=6810;
					out<=10;
				end
				if(in == 3) begin
					state<=1476;
					out<=11;
				end
				if(in == 4) begin
					state<=5365;
					out<=12;
				end
			end
			2921: begin
				if(in == 0) begin
					state<=2922;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=6811;
					out<=15;
				end
				if(in == 3) begin
					state<=1477;
					out<=16;
				end
				if(in == 4) begin
					state<=5366;
					out<=17;
				end
			end
			2922: begin
				if(in == 0) begin
					state<=2923;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=6812;
					out<=20;
				end
				if(in == 3) begin
					state<=1478;
					out<=21;
				end
				if(in == 4) begin
					state<=5367;
					out<=22;
				end
			end
			2923: begin
				if(in == 0) begin
					state<=2924;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=6813;
					out<=25;
				end
				if(in == 3) begin
					state<=1479;
					out<=26;
				end
				if(in == 4) begin
					state<=5368;
					out<=27;
				end
			end
			2924: begin
				if(in == 0) begin
					state<=2925;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=6814;
					out<=30;
				end
				if(in == 3) begin
					state<=1480;
					out<=31;
				end
				if(in == 4) begin
					state<=5369;
					out<=32;
				end
			end
			2925: begin
				if(in == 0) begin
					state<=2926;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=6815;
					out<=35;
				end
				if(in == 3) begin
					state<=1481;
					out<=36;
				end
				if(in == 4) begin
					state<=5370;
					out<=37;
				end
			end
			2926: begin
				if(in == 0) begin
					state<=2927;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=6816;
					out<=40;
				end
				if(in == 3) begin
					state<=1482;
					out<=41;
				end
				if(in == 4) begin
					state<=5371;
					out<=42;
				end
			end
			2927: begin
				if(in == 0) begin
					state<=2928;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=6817;
					out<=45;
				end
				if(in == 3) begin
					state<=1483;
					out<=46;
				end
				if(in == 4) begin
					state<=5372;
					out<=47;
				end
			end
			2928: begin
				if(in == 0) begin
					state<=2325;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=6214;
					out<=50;
				end
				if(in == 3) begin
					state<=327;
					out<=51;
				end
				if(in == 4) begin
					state<=4225;
					out<=52;
				end
			end
			2929: begin
				if(in == 0) begin
					state<=2930;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=6819;
					out<=55;
				end
				if(in == 3) begin
					state<=347;
					out<=56;
				end
				if(in == 4) begin
					state<=4245;
					out<=57;
				end
			end
			2930: begin
				if(in == 0) begin
					state<=2931;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=6820;
					out<=60;
				end
				if(in == 3) begin
					state<=348;
					out<=61;
				end
				if(in == 4) begin
					state<=4246;
					out<=62;
				end
			end
			2931: begin
				if(in == 0) begin
					state<=2932;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=6821;
					out<=65;
				end
				if(in == 3) begin
					state<=349;
					out<=66;
				end
				if(in == 4) begin
					state<=4247;
					out<=67;
				end
			end
			2932: begin
				if(in == 0) begin
					state<=2933;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=6822;
					out<=70;
				end
				if(in == 3) begin
					state<=350;
					out<=71;
				end
				if(in == 4) begin
					state<=4248;
					out<=72;
				end
			end
			2933: begin
				if(in == 0) begin
					state<=2934;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=6823;
					out<=75;
				end
				if(in == 3) begin
					state<=351;
					out<=76;
				end
				if(in == 4) begin
					state<=4249;
					out<=77;
				end
			end
			2934: begin
				if(in == 0) begin
					state<=2935;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=6824;
					out<=80;
				end
				if(in == 3) begin
					state<=352;
					out<=81;
				end
				if(in == 4) begin
					state<=4250;
					out<=82;
				end
			end
			2935: begin
				if(in == 0) begin
					state<=2936;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=6825;
					out<=85;
				end
				if(in == 3) begin
					state<=353;
					out<=86;
				end
				if(in == 4) begin
					state<=4251;
					out<=87;
				end
			end
			2936: begin
				if(in == 0) begin
					state<=2937;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=6826;
					out<=90;
				end
				if(in == 3) begin
					state<=354;
					out<=91;
				end
				if(in == 4) begin
					state<=4252;
					out<=92;
				end
			end
			2937: begin
				if(in == 0) begin
					state<=2938;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=6827;
					out<=95;
				end
				if(in == 3) begin
					state<=355;
					out<=96;
				end
				if(in == 4) begin
					state<=4253;
					out<=97;
				end
			end
			2938: begin
				if(in == 0) begin
					state<=2939;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=6828;
					out<=100;
				end
				if(in == 3) begin
					state<=356;
					out<=101;
				end
				if(in == 4) begin
					state<=4254;
					out<=102;
				end
			end
			2939: begin
				if(in == 0) begin
					state<=2940;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=6829;
					out<=105;
				end
				if(in == 3) begin
					state<=357;
					out<=106;
				end
				if(in == 4) begin
					state<=4255;
					out<=107;
				end
			end
			2940: begin
				if(in == 0) begin
					state<=2941;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=6830;
					out<=110;
				end
				if(in == 3) begin
					state<=358;
					out<=111;
				end
				if(in == 4) begin
					state<=4256;
					out<=112;
				end
			end
			2941: begin
				if(in == 0) begin
					state<=2942;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=6831;
					out<=115;
				end
				if(in == 3) begin
					state<=359;
					out<=116;
				end
				if(in == 4) begin
					state<=4257;
					out<=117;
				end
			end
			2942: begin
				if(in == 0) begin
					state<=2943;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=6832;
					out<=120;
				end
				if(in == 3) begin
					state<=360;
					out<=121;
				end
				if(in == 4) begin
					state<=4258;
					out<=122;
				end
			end
			2943: begin
				if(in == 0) begin
					state<=2944;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=6833;
					out<=125;
				end
				if(in == 3) begin
					state<=361;
					out<=126;
				end
				if(in == 4) begin
					state<=4259;
					out<=127;
				end
			end
			2944: begin
				if(in == 0) begin
					state<=2945;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=6834;
					out<=130;
				end
				if(in == 3) begin
					state<=362;
					out<=131;
				end
				if(in == 4) begin
					state<=4260;
					out<=132;
				end
			end
			2945: begin
				if(in == 0) begin
					state<=2946;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=6835;
					out<=135;
				end
				if(in == 3) begin
					state<=363;
					out<=136;
				end
				if(in == 4) begin
					state<=4261;
					out<=137;
				end
			end
			2946: begin
				if(in == 0) begin
					state<=2947;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=6836;
					out<=140;
				end
				if(in == 3) begin
					state<=364;
					out<=141;
				end
				if(in == 4) begin
					state<=4262;
					out<=142;
				end
			end
			2947: begin
				if(in == 0) begin
					state<=2948;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=6837;
					out<=145;
				end
				if(in == 3) begin
					state<=365;
					out<=146;
				end
				if(in == 4) begin
					state<=4263;
					out<=147;
				end
			end
			2948: begin
				if(in == 0) begin
					state<=2949;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=6838;
					out<=150;
				end
				if(in == 3) begin
					state<=366;
					out<=151;
				end
				if(in == 4) begin
					state<=4264;
					out<=152;
				end
			end
			2949: begin
				if(in == 0) begin
					state<=2950;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=6839;
					out<=155;
				end
				if(in == 3) begin
					state<=367;
					out<=156;
				end
				if(in == 4) begin
					state<=4265;
					out<=157;
				end
			end
			2950: begin
				if(in == 0) begin
					state<=2951;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=6840;
					out<=160;
				end
				if(in == 3) begin
					state<=368;
					out<=161;
				end
				if(in == 4) begin
					state<=4266;
					out<=162;
				end
			end
			2951: begin
				if(in == 0) begin
					state<=2952;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=6841;
					out<=165;
				end
				if(in == 3) begin
					state<=369;
					out<=166;
				end
				if(in == 4) begin
					state<=4267;
					out<=167;
				end
			end
			2952: begin
				if(in == 0) begin
					state<=2953;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=6842;
					out<=170;
				end
				if(in == 3) begin
					state<=370;
					out<=171;
				end
				if(in == 4) begin
					state<=4268;
					out<=172;
				end
			end
			2953: begin
				if(in == 0) begin
					state<=2954;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=6843;
					out<=175;
				end
				if(in == 3) begin
					state<=371;
					out<=176;
				end
				if(in == 4) begin
					state<=4269;
					out<=177;
				end
			end
			2954: begin
				if(in == 0) begin
					state<=2955;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=6844;
					out<=180;
				end
				if(in == 3) begin
					state<=372;
					out<=181;
				end
				if(in == 4) begin
					state<=4270;
					out<=182;
				end
			end
			2955: begin
				if(in == 0) begin
					state<=2956;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=6845;
					out<=185;
				end
				if(in == 3) begin
					state<=373;
					out<=186;
				end
				if(in == 4) begin
					state<=4271;
					out<=187;
				end
			end
			2956: begin
				if(in == 0) begin
					state<=2957;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=6846;
					out<=190;
				end
				if(in == 3) begin
					state<=374;
					out<=191;
				end
				if(in == 4) begin
					state<=4272;
					out<=192;
				end
			end
			2957: begin
				if(in == 0) begin
					state<=2958;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=6847;
					out<=195;
				end
				if(in == 3) begin
					state<=375;
					out<=196;
				end
				if(in == 4) begin
					state<=4273;
					out<=197;
				end
			end
			2958: begin
				if(in == 0) begin
					state<=2959;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=6848;
					out<=200;
				end
				if(in == 3) begin
					state<=376;
					out<=201;
				end
				if(in == 4) begin
					state<=4274;
					out<=202;
				end
			end
			2959: begin
				if(in == 0) begin
					state<=2960;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=6849;
					out<=205;
				end
				if(in == 3) begin
					state<=377;
					out<=206;
				end
				if(in == 4) begin
					state<=4275;
					out<=207;
				end
			end
			2960: begin
				if(in == 0) begin
					state<=2961;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=6850;
					out<=210;
				end
				if(in == 3) begin
					state<=378;
					out<=211;
				end
				if(in == 4) begin
					state<=4276;
					out<=212;
				end
			end
			2961: begin
				if(in == 0) begin
					state<=2962;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=6851;
					out<=215;
				end
				if(in == 3) begin
					state<=379;
					out<=216;
				end
				if(in == 4) begin
					state<=4277;
					out<=217;
				end
			end
			2962: begin
				if(in == 0) begin
					state<=2963;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=6852;
					out<=220;
				end
				if(in == 3) begin
					state<=380;
					out<=221;
				end
				if(in == 4) begin
					state<=4278;
					out<=222;
				end
			end
			2963: begin
				if(in == 0) begin
					state<=2964;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=6853;
					out<=225;
				end
				if(in == 3) begin
					state<=381;
					out<=226;
				end
				if(in == 4) begin
					state<=4279;
					out<=227;
				end
			end
			2964: begin
				if(in == 0) begin
					state<=2965;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=6854;
					out<=230;
				end
				if(in == 3) begin
					state<=382;
					out<=231;
				end
				if(in == 4) begin
					state<=4280;
					out<=232;
				end
			end
			2965: begin
				if(in == 0) begin
					state<=2966;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=6855;
					out<=235;
				end
				if(in == 3) begin
					state<=383;
					out<=236;
				end
				if(in == 4) begin
					state<=4281;
					out<=237;
				end
			end
			2966: begin
				if(in == 0) begin
					state<=2967;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=6856;
					out<=240;
				end
				if(in == 3) begin
					state<=384;
					out<=241;
				end
				if(in == 4) begin
					state<=4282;
					out<=242;
				end
			end
			2967: begin
				if(in == 0) begin
					state<=2968;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=6857;
					out<=245;
				end
				if(in == 3) begin
					state<=385;
					out<=246;
				end
				if(in == 4) begin
					state<=4283;
					out<=247;
				end
			end
			2968: begin
				if(in == 0) begin
					state<=2969;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=6858;
					out<=250;
				end
				if(in == 3) begin
					state<=386;
					out<=251;
				end
				if(in == 4) begin
					state<=4284;
					out<=252;
				end
			end
			2969: begin
				if(in == 0) begin
					state<=2970;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=6859;
					out<=255;
				end
				if(in == 3) begin
					state<=387;
					out<=0;
				end
				if(in == 4) begin
					state<=4285;
					out<=1;
				end
			end
			2970: begin
				if(in == 0) begin
					state<=2971;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=6860;
					out<=4;
				end
				if(in == 3) begin
					state<=388;
					out<=5;
				end
				if(in == 4) begin
					state<=4286;
					out<=6;
				end
			end
			2971: begin
				if(in == 0) begin
					state<=2972;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=6861;
					out<=9;
				end
				if(in == 3) begin
					state<=389;
					out<=10;
				end
				if(in == 4) begin
					state<=4287;
					out<=11;
				end
			end
			2972: begin
				if(in == 0) begin
					state<=2973;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=6862;
					out<=14;
				end
				if(in == 3) begin
					state<=390;
					out<=15;
				end
				if(in == 4) begin
					state<=4288;
					out<=16;
				end
			end
			2973: begin
				if(in == 0) begin
					state<=2974;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=6863;
					out<=19;
				end
				if(in == 3) begin
					state<=391;
					out<=20;
				end
				if(in == 4) begin
					state<=4289;
					out<=21;
				end
			end
			2974: begin
				if(in == 0) begin
					state<=2975;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=6864;
					out<=24;
				end
				if(in == 3) begin
					state<=392;
					out<=25;
				end
				if(in == 4) begin
					state<=4290;
					out<=26;
				end
			end
			2975: begin
				if(in == 0) begin
					state<=2976;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=6865;
					out<=29;
				end
				if(in == 3) begin
					state<=393;
					out<=30;
				end
				if(in == 4) begin
					state<=4291;
					out<=31;
				end
			end
			2976: begin
				if(in == 0) begin
					state<=2977;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=6866;
					out<=34;
				end
				if(in == 3) begin
					state<=394;
					out<=35;
				end
				if(in == 4) begin
					state<=4292;
					out<=36;
				end
			end
			2977: begin
				if(in == 0) begin
					state<=2978;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=6867;
					out<=39;
				end
				if(in == 3) begin
					state<=395;
					out<=40;
				end
				if(in == 4) begin
					state<=4293;
					out<=41;
				end
			end
			2978: begin
				if(in == 0) begin
					state<=2979;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=6868;
					out<=44;
				end
				if(in == 3) begin
					state<=999;
					out<=45;
				end
				if(in == 4) begin
					state<=4897;
					out<=46;
				end
			end
			2979: begin
				if(in == 0) begin
					state<=2980;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=6869;
					out<=49;
				end
				if(in == 3) begin
					state<=1000;
					out<=50;
				end
				if(in == 4) begin
					state<=4898;
					out<=51;
				end
			end
			2980: begin
				if(in == 0) begin
					state<=2981;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=6870;
					out<=54;
				end
				if(in == 3) begin
					state<=1001;
					out<=55;
				end
				if(in == 4) begin
					state<=4899;
					out<=56;
				end
			end
			2981: begin
				if(in == 0) begin
					state<=2982;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=6871;
					out<=59;
				end
				if(in == 3) begin
					state<=1002;
					out<=60;
				end
				if(in == 4) begin
					state<=4900;
					out<=61;
				end
			end
			2982: begin
				if(in == 0) begin
					state<=2983;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=6872;
					out<=64;
				end
				if(in == 3) begin
					state<=1003;
					out<=65;
				end
				if(in == 4) begin
					state<=4901;
					out<=66;
				end
			end
			2983: begin
				if(in == 0) begin
					state<=2984;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=6873;
					out<=69;
				end
				if(in == 3) begin
					state<=1004;
					out<=70;
				end
				if(in == 4) begin
					state<=4902;
					out<=71;
				end
			end
			2984: begin
				if(in == 0) begin
					state<=2985;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=6874;
					out<=74;
				end
				if(in == 3) begin
					state<=1005;
					out<=75;
				end
				if(in == 4) begin
					state<=4903;
					out<=76;
				end
			end
			2985: begin
				if(in == 0) begin
					state<=2986;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=6875;
					out<=79;
				end
				if(in == 3) begin
					state<=1006;
					out<=80;
				end
				if(in == 4) begin
					state<=4904;
					out<=81;
				end
			end
			2986: begin
				if(in == 0) begin
					state<=2987;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=6876;
					out<=84;
				end
				if(in == 3) begin
					state<=1007;
					out<=85;
				end
				if(in == 4) begin
					state<=4905;
					out<=86;
				end
			end
			2987: begin
				if(in == 0) begin
					state<=2988;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=6877;
					out<=89;
				end
				if(in == 3) begin
					state<=1008;
					out<=90;
				end
				if(in == 4) begin
					state<=4906;
					out<=91;
				end
			end
			2988: begin
				if(in == 0) begin
					state<=2989;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=6878;
					out<=94;
				end
				if(in == 3) begin
					state<=1009;
					out<=95;
				end
				if(in == 4) begin
					state<=4907;
					out<=96;
				end
			end
			2989: begin
				if(in == 0) begin
					state<=2990;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=6879;
					out<=99;
				end
				if(in == 3) begin
					state<=1010;
					out<=100;
				end
				if(in == 4) begin
					state<=4908;
					out<=101;
				end
			end
			2990: begin
				if(in == 0) begin
					state<=2991;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=6880;
					out<=104;
				end
				if(in == 3) begin
					state<=1011;
					out<=105;
				end
				if(in == 4) begin
					state<=4909;
					out<=106;
				end
			end
			2991: begin
				if(in == 0) begin
					state<=2992;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=6881;
					out<=109;
				end
				if(in == 3) begin
					state<=1012;
					out<=110;
				end
				if(in == 4) begin
					state<=4910;
					out<=111;
				end
			end
			2992: begin
				if(in == 0) begin
					state<=2993;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=6882;
					out<=114;
				end
				if(in == 3) begin
					state<=1013;
					out<=115;
				end
				if(in == 4) begin
					state<=4911;
					out<=116;
				end
			end
			2993: begin
				if(in == 0) begin
					state<=2994;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=6883;
					out<=119;
				end
				if(in == 3) begin
					state<=1014;
					out<=120;
				end
				if(in == 4) begin
					state<=4912;
					out<=121;
				end
			end
			2994: begin
				if(in == 0) begin
					state<=2995;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=6884;
					out<=124;
				end
				if(in == 3) begin
					state<=1015;
					out<=125;
				end
				if(in == 4) begin
					state<=4913;
					out<=126;
				end
			end
			2995: begin
				if(in == 0) begin
					state<=2996;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=6885;
					out<=129;
				end
				if(in == 3) begin
					state<=1016;
					out<=130;
				end
				if(in == 4) begin
					state<=4914;
					out<=131;
				end
			end
			2996: begin
				if(in == 0) begin
					state<=2997;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=6886;
					out<=134;
				end
				if(in == 3) begin
					state<=1017;
					out<=135;
				end
				if(in == 4) begin
					state<=4915;
					out<=136;
				end
			end
			2997: begin
				if(in == 0) begin
					state<=2998;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=6887;
					out<=139;
				end
				if(in == 3) begin
					state<=1018;
					out<=140;
				end
				if(in == 4) begin
					state<=4916;
					out<=141;
				end
			end
			2998: begin
				if(in == 0) begin
					state<=2999;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=6888;
					out<=144;
				end
				if(in == 3) begin
					state<=1019;
					out<=145;
				end
				if(in == 4) begin
					state<=4917;
					out<=146;
				end
			end
			2999: begin
				if(in == 0) begin
					state<=3000;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=6889;
					out<=149;
				end
				if(in == 3) begin
					state<=1020;
					out<=150;
				end
				if(in == 4) begin
					state<=4918;
					out<=151;
				end
			end
			3000: begin
				if(in == 0) begin
					state<=3001;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=6890;
					out<=154;
				end
				if(in == 3) begin
					state<=1021;
					out<=155;
				end
				if(in == 4) begin
					state<=4919;
					out<=156;
				end
			end
			3001: begin
				if(in == 0) begin
					state<=3002;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=6891;
					out<=159;
				end
				if(in == 3) begin
					state<=1022;
					out<=160;
				end
				if(in == 4) begin
					state<=4920;
					out<=161;
				end
			end
			3002: begin
				if(in == 0) begin
					state<=3003;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=6892;
					out<=164;
				end
				if(in == 3) begin
					state<=1023;
					out<=165;
				end
				if(in == 4) begin
					state<=4921;
					out<=166;
				end
			end
			3003: begin
				if(in == 0) begin
					state<=3004;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=6893;
					out<=169;
				end
				if(in == 3) begin
					state<=1024;
					out<=170;
				end
				if(in == 4) begin
					state<=4922;
					out<=171;
				end
			end
			3004: begin
				if(in == 0) begin
					state<=3005;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=6894;
					out<=174;
				end
				if(in == 3) begin
					state<=1025;
					out<=175;
				end
				if(in == 4) begin
					state<=4923;
					out<=176;
				end
			end
			3005: begin
				if(in == 0) begin
					state<=3006;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=6895;
					out<=179;
				end
				if(in == 3) begin
					state<=1026;
					out<=180;
				end
				if(in == 4) begin
					state<=4924;
					out<=181;
				end
			end
			3006: begin
				if(in == 0) begin
					state<=3007;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=6896;
					out<=184;
				end
				if(in == 3) begin
					state<=1027;
					out<=185;
				end
				if(in == 4) begin
					state<=4925;
					out<=186;
				end
			end
			3007: begin
				if(in == 0) begin
					state<=3008;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=6897;
					out<=189;
				end
				if(in == 3) begin
					state<=1028;
					out<=190;
				end
				if(in == 4) begin
					state<=4926;
					out<=191;
				end
			end
			3008: begin
				if(in == 0) begin
					state<=3009;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=6898;
					out<=194;
				end
				if(in == 3) begin
					state<=1029;
					out<=195;
				end
				if(in == 4) begin
					state<=4927;
					out<=196;
				end
			end
			3009: begin
				if(in == 0) begin
					state<=3010;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=6899;
					out<=199;
				end
				if(in == 3) begin
					state<=396;
					out<=200;
				end
				if(in == 4) begin
					state<=4294;
					out<=201;
				end
			end
			3010: begin
				if(in == 0) begin
					state<=3011;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=6900;
					out<=204;
				end
				if(in == 3) begin
					state<=397;
					out<=205;
				end
				if(in == 4) begin
					state<=4295;
					out<=206;
				end
			end
			3011: begin
				if(in == 0) begin
					state<=3012;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=6901;
					out<=209;
				end
				if(in == 3) begin
					state<=398;
					out<=210;
				end
				if(in == 4) begin
					state<=4296;
					out<=211;
				end
			end
			3012: begin
				if(in == 0) begin
					state<=3013;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=6902;
					out<=214;
				end
				if(in == 3) begin
					state<=399;
					out<=215;
				end
				if(in == 4) begin
					state<=4297;
					out<=216;
				end
			end
			3013: begin
				if(in == 0) begin
					state<=3014;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=6903;
					out<=219;
				end
				if(in == 3) begin
					state<=400;
					out<=220;
				end
				if(in == 4) begin
					state<=4298;
					out<=221;
				end
			end
			3014: begin
				if(in == 0) begin
					state<=3015;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=6904;
					out<=224;
				end
				if(in == 3) begin
					state<=401;
					out<=225;
				end
				if(in == 4) begin
					state<=4299;
					out<=226;
				end
			end
			3015: begin
				if(in == 0) begin
					state<=3016;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=6905;
					out<=229;
				end
				if(in == 3) begin
					state<=402;
					out<=230;
				end
				if(in == 4) begin
					state<=4300;
					out<=231;
				end
			end
			3016: begin
				if(in == 0) begin
					state<=3017;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=6906;
					out<=234;
				end
				if(in == 3) begin
					state<=403;
					out<=235;
				end
				if(in == 4) begin
					state<=4301;
					out<=236;
				end
			end
			3017: begin
				if(in == 0) begin
					state<=3018;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=6907;
					out<=239;
				end
				if(in == 3) begin
					state<=404;
					out<=240;
				end
				if(in == 4) begin
					state<=4302;
					out<=241;
				end
			end
			3018: begin
				if(in == 0) begin
					state<=3019;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=6908;
					out<=244;
				end
				if(in == 3) begin
					state<=405;
					out<=245;
				end
				if(in == 4) begin
					state<=4303;
					out<=246;
				end
			end
			3019: begin
				if(in == 0) begin
					state<=3020;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=6909;
					out<=249;
				end
				if(in == 3) begin
					state<=406;
					out<=250;
				end
				if(in == 4) begin
					state<=4304;
					out<=251;
				end
			end
			3020: begin
				if(in == 0) begin
					state<=3021;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=6910;
					out<=254;
				end
				if(in == 3) begin
					state<=407;
					out<=255;
				end
				if(in == 4) begin
					state<=4305;
					out<=0;
				end
			end
			3021: begin
				if(in == 0) begin
					state<=3022;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=6911;
					out<=3;
				end
				if(in == 3) begin
					state<=408;
					out<=4;
				end
				if(in == 4) begin
					state<=4306;
					out<=5;
				end
			end
			3022: begin
				if(in == 0) begin
					state<=3023;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=6912;
					out<=8;
				end
				if(in == 3) begin
					state<=409;
					out<=9;
				end
				if(in == 4) begin
					state<=4307;
					out<=10;
				end
			end
			3023: begin
				if(in == 0) begin
					state<=3024;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=6913;
					out<=13;
				end
				if(in == 3) begin
					state<=410;
					out<=14;
				end
				if(in == 4) begin
					state<=4308;
					out<=15;
				end
			end
			3024: begin
				if(in == 0) begin
					state<=3025;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=6914;
					out<=18;
				end
				if(in == 3) begin
					state<=411;
					out<=19;
				end
				if(in == 4) begin
					state<=4309;
					out<=20;
				end
			end
			3025: begin
				if(in == 0) begin
					state<=3026;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=6915;
					out<=23;
				end
				if(in == 3) begin
					state<=412;
					out<=24;
				end
				if(in == 4) begin
					state<=4310;
					out<=25;
				end
			end
			3026: begin
				if(in == 0) begin
					state<=3027;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=6916;
					out<=28;
				end
				if(in == 3) begin
					state<=413;
					out<=29;
				end
				if(in == 4) begin
					state<=4311;
					out<=30;
				end
			end
			3027: begin
				if(in == 0) begin
					state<=3028;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=6917;
					out<=33;
				end
				if(in == 3) begin
					state<=414;
					out<=34;
				end
				if(in == 4) begin
					state<=4312;
					out<=35;
				end
			end
			3028: begin
				if(in == 0) begin
					state<=3029;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=6918;
					out<=38;
				end
				if(in == 3) begin
					state<=1030;
					out<=39;
				end
				if(in == 4) begin
					state<=4928;
					out<=40;
				end
			end
			3029: begin
				if(in == 0) begin
					state<=3030;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=6919;
					out<=43;
				end
				if(in == 3) begin
					state<=1031;
					out<=44;
				end
				if(in == 4) begin
					state<=4929;
					out<=45;
				end
			end
			3030: begin
				if(in == 0) begin
					state<=3031;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=6920;
					out<=48;
				end
				if(in == 3) begin
					state<=1032;
					out<=49;
				end
				if(in == 4) begin
					state<=4930;
					out<=50;
				end
			end
			3031: begin
				if(in == 0) begin
					state<=3032;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=6921;
					out<=53;
				end
				if(in == 3) begin
					state<=1033;
					out<=54;
				end
				if(in == 4) begin
					state<=4931;
					out<=55;
				end
			end
			3032: begin
				if(in == 0) begin
					state<=3033;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=6922;
					out<=58;
				end
				if(in == 3) begin
					state<=1034;
					out<=59;
				end
				if(in == 4) begin
					state<=4932;
					out<=60;
				end
			end
			3033: begin
				if(in == 0) begin
					state<=3034;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=6923;
					out<=63;
				end
				if(in == 3) begin
					state<=1035;
					out<=64;
				end
				if(in == 4) begin
					state<=4933;
					out<=65;
				end
			end
			3034: begin
				if(in == 0) begin
					state<=3035;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=6924;
					out<=68;
				end
				if(in == 3) begin
					state<=1036;
					out<=69;
				end
				if(in == 4) begin
					state<=4934;
					out<=70;
				end
			end
			3035: begin
				if(in == 0) begin
					state<=3036;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=6925;
					out<=73;
				end
				if(in == 3) begin
					state<=1037;
					out<=74;
				end
				if(in == 4) begin
					state<=4935;
					out<=75;
				end
			end
			3036: begin
				if(in == 0) begin
					state<=3037;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=6926;
					out<=78;
				end
				if(in == 3) begin
					state<=1038;
					out<=79;
				end
				if(in == 4) begin
					state<=4936;
					out<=80;
				end
			end
			3037: begin
				if(in == 0) begin
					state<=3038;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=6927;
					out<=83;
				end
				if(in == 3) begin
					state<=1039;
					out<=84;
				end
				if(in == 4) begin
					state<=4937;
					out<=85;
				end
			end
			3038: begin
				if(in == 0) begin
					state<=3039;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=6928;
					out<=88;
				end
				if(in == 3) begin
					state<=1040;
					out<=89;
				end
				if(in == 4) begin
					state<=4938;
					out<=90;
				end
			end
			3039: begin
				if(in == 0) begin
					state<=3040;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=6929;
					out<=93;
				end
				if(in == 3) begin
					state<=1041;
					out<=94;
				end
				if(in == 4) begin
					state<=4939;
					out<=95;
				end
			end
			3040: begin
				if(in == 0) begin
					state<=3041;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=6930;
					out<=98;
				end
				if(in == 3) begin
					state<=1042;
					out<=99;
				end
				if(in == 4) begin
					state<=4940;
					out<=100;
				end
			end
			3041: begin
				if(in == 0) begin
					state<=3042;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=6931;
					out<=103;
				end
				if(in == 3) begin
					state<=1043;
					out<=104;
				end
				if(in == 4) begin
					state<=4941;
					out<=105;
				end
			end
			3042: begin
				if(in == 0) begin
					state<=3043;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=6932;
					out<=108;
				end
				if(in == 3) begin
					state<=1044;
					out<=109;
				end
				if(in == 4) begin
					state<=4942;
					out<=110;
				end
			end
			3043: begin
				if(in == 0) begin
					state<=3044;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=6933;
					out<=113;
				end
				if(in == 3) begin
					state<=1045;
					out<=114;
				end
				if(in == 4) begin
					state<=4943;
					out<=115;
				end
			end
			3044: begin
				if(in == 0) begin
					state<=3045;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=6934;
					out<=118;
				end
				if(in == 3) begin
					state<=1046;
					out<=119;
				end
				if(in == 4) begin
					state<=4944;
					out<=120;
				end
			end
			3045: begin
				if(in == 0) begin
					state<=3046;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=6935;
					out<=123;
				end
				if(in == 3) begin
					state<=1047;
					out<=124;
				end
				if(in == 4) begin
					state<=4945;
					out<=125;
				end
			end
			3046: begin
				if(in == 0) begin
					state<=3047;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=6936;
					out<=128;
				end
				if(in == 3) begin
					state<=1048;
					out<=129;
				end
				if(in == 4) begin
					state<=4946;
					out<=130;
				end
			end
			3047: begin
				if(in == 0) begin
					state<=3048;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=6937;
					out<=133;
				end
				if(in == 3) begin
					state<=1049;
					out<=134;
				end
				if(in == 4) begin
					state<=4947;
					out<=135;
				end
			end
			3048: begin
				if(in == 0) begin
					state<=3049;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=6938;
					out<=138;
				end
				if(in == 3) begin
					state<=1050;
					out<=139;
				end
				if(in == 4) begin
					state<=4948;
					out<=140;
				end
			end
			3049: begin
				if(in == 0) begin
					state<=3050;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=6939;
					out<=143;
				end
				if(in == 3) begin
					state<=1051;
					out<=144;
				end
				if(in == 4) begin
					state<=4949;
					out<=145;
				end
			end
			3050: begin
				if(in == 0) begin
					state<=3051;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=6940;
					out<=148;
				end
				if(in == 3) begin
					state<=1052;
					out<=149;
				end
				if(in == 4) begin
					state<=4950;
					out<=150;
				end
			end
			3051: begin
				if(in == 0) begin
					state<=3052;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=6941;
					out<=153;
				end
				if(in == 3) begin
					state<=1053;
					out<=154;
				end
				if(in == 4) begin
					state<=4951;
					out<=155;
				end
			end
			3052: begin
				if(in == 0) begin
					state<=3053;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=6942;
					out<=158;
				end
				if(in == 3) begin
					state<=1054;
					out<=159;
				end
				if(in == 4) begin
					state<=4952;
					out<=160;
				end
			end
			3053: begin
				if(in == 0) begin
					state<=3054;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=6943;
					out<=163;
				end
				if(in == 3) begin
					state<=1055;
					out<=164;
				end
				if(in == 4) begin
					state<=4953;
					out<=165;
				end
			end
			3054: begin
				if(in == 0) begin
					state<=3055;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=6944;
					out<=168;
				end
				if(in == 3) begin
					state<=1056;
					out<=169;
				end
				if(in == 4) begin
					state<=4954;
					out<=170;
				end
			end
			3055: begin
				if(in == 0) begin
					state<=3056;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=6945;
					out<=173;
				end
				if(in == 3) begin
					state<=1057;
					out<=174;
				end
				if(in == 4) begin
					state<=4955;
					out<=175;
				end
			end
			3056: begin
				if(in == 0) begin
					state<=3057;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=6946;
					out<=178;
				end
				if(in == 3) begin
					state<=1058;
					out<=179;
				end
				if(in == 4) begin
					state<=4956;
					out<=180;
				end
			end
			3057: begin
				if(in == 0) begin
					state<=3058;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=6947;
					out<=183;
				end
				if(in == 3) begin
					state<=1059;
					out<=184;
				end
				if(in == 4) begin
					state<=4957;
					out<=185;
				end
			end
			3058: begin
				if(in == 0) begin
					state<=3059;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=6948;
					out<=188;
				end
				if(in == 3) begin
					state<=1060;
					out<=189;
				end
				if(in == 4) begin
					state<=4958;
					out<=190;
				end
			end
			3059: begin
				if(in == 0) begin
					state<=3060;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=6949;
					out<=193;
				end
				if(in == 3) begin
					state<=1061;
					out<=194;
				end
				if(in == 4) begin
					state<=4959;
					out<=195;
				end
			end
			3060: begin
				if(in == 0) begin
					state<=3061;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=6950;
					out<=198;
				end
				if(in == 3) begin
					state<=1062;
					out<=199;
				end
				if(in == 4) begin
					state<=4960;
					out<=200;
				end
			end
			3061: begin
				if(in == 0) begin
					state<=3062;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=6951;
					out<=203;
				end
				if(in == 3) begin
					state<=1063;
					out<=204;
				end
				if(in == 4) begin
					state<=4961;
					out<=205;
				end
			end
			3062: begin
				if(in == 0) begin
					state<=3063;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=6952;
					out<=208;
				end
				if(in == 3) begin
					state<=1064;
					out<=209;
				end
				if(in == 4) begin
					state<=4962;
					out<=210;
				end
			end
			3063: begin
				if(in == 0) begin
					state<=3064;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=6953;
					out<=213;
				end
				if(in == 3) begin
					state<=1065;
					out<=214;
				end
				if(in == 4) begin
					state<=4963;
					out<=215;
				end
			end
			3064: begin
				if(in == 0) begin
					state<=3065;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=6954;
					out<=218;
				end
				if(in == 3) begin
					state<=1066;
					out<=219;
				end
				if(in == 4) begin
					state<=4964;
					out<=220;
				end
			end
			3065: begin
				if(in == 0) begin
					state<=3066;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=6955;
					out<=223;
				end
				if(in == 3) begin
					state<=1067;
					out<=224;
				end
				if(in == 4) begin
					state<=4965;
					out<=225;
				end
			end
			3066: begin
				if(in == 0) begin
					state<=3067;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=6956;
					out<=228;
				end
				if(in == 3) begin
					state<=1068;
					out<=229;
				end
				if(in == 4) begin
					state<=4966;
					out<=230;
				end
			end
			3067: begin
				if(in == 0) begin
					state<=3068;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=6957;
					out<=233;
				end
				if(in == 3) begin
					state<=1069;
					out<=234;
				end
				if(in == 4) begin
					state<=4967;
					out<=235;
				end
			end
			3068: begin
				if(in == 0) begin
					state<=3069;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=6958;
					out<=238;
				end
				if(in == 3) begin
					state<=1070;
					out<=239;
				end
				if(in == 4) begin
					state<=4968;
					out<=240;
				end
			end
			3069: begin
				if(in == 0) begin
					state<=3070;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=6959;
					out<=243;
				end
				if(in == 3) begin
					state<=1071;
					out<=244;
				end
				if(in == 4) begin
					state<=4969;
					out<=245;
				end
			end
			3070: begin
				if(in == 0) begin
					state<=3071;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=6960;
					out<=248;
				end
				if(in == 3) begin
					state<=1072;
					out<=249;
				end
				if(in == 4) begin
					state<=4970;
					out<=250;
				end
			end
			3071: begin
				if(in == 0) begin
					state<=3072;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=6961;
					out<=253;
				end
				if(in == 3) begin
					state<=1073;
					out<=254;
				end
				if(in == 4) begin
					state<=4971;
					out<=255;
				end
			end
			3072: begin
				if(in == 0) begin
					state<=3073;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=6962;
					out<=2;
				end
				if(in == 3) begin
					state<=1074;
					out<=3;
				end
				if(in == 4) begin
					state<=4972;
					out<=4;
				end
			end
			3073: begin
				if(in == 0) begin
					state<=3074;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=6963;
					out<=7;
				end
				if(in == 3) begin
					state<=1075;
					out<=8;
				end
				if(in == 4) begin
					state<=4973;
					out<=9;
				end
			end
			3074: begin
				if(in == 0) begin
					state<=3075;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=6964;
					out<=12;
				end
				if(in == 3) begin
					state<=1076;
					out<=13;
				end
				if(in == 4) begin
					state<=4974;
					out<=14;
				end
			end
			3075: begin
				if(in == 0) begin
					state<=3076;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=6965;
					out<=17;
				end
				if(in == 3) begin
					state<=1077;
					out<=18;
				end
				if(in == 4) begin
					state<=4975;
					out<=19;
				end
			end
			3076: begin
				if(in == 0) begin
					state<=3077;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=6966;
					out<=22;
				end
				if(in == 3) begin
					state<=1078;
					out<=23;
				end
				if(in == 4) begin
					state<=4976;
					out<=24;
				end
			end
			3077: begin
				if(in == 0) begin
					state<=3078;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=6967;
					out<=27;
				end
				if(in == 3) begin
					state<=1079;
					out<=28;
				end
				if(in == 4) begin
					state<=4977;
					out<=29;
				end
			end
			3078: begin
				if(in == 0) begin
					state<=3079;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=6968;
					out<=32;
				end
				if(in == 3) begin
					state<=1080;
					out<=33;
				end
				if(in == 4) begin
					state<=4978;
					out<=34;
				end
			end
			3079: begin
				if(in == 0) begin
					state<=3080;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=6969;
					out<=37;
				end
				if(in == 3) begin
					state<=1081;
					out<=38;
				end
				if(in == 4) begin
					state<=4979;
					out<=39;
				end
			end
			3080: begin
				if(in == 0) begin
					state<=3081;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=6970;
					out<=42;
				end
				if(in == 3) begin
					state<=1082;
					out<=43;
				end
				if(in == 4) begin
					state<=4980;
					out<=44;
				end
			end
			3081: begin
				if(in == 0) begin
					state<=3082;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=6971;
					out<=47;
				end
				if(in == 3) begin
					state<=1083;
					out<=48;
				end
				if(in == 4) begin
					state<=4981;
					out<=49;
				end
			end
			3082: begin
				if(in == 0) begin
					state<=3083;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=6972;
					out<=52;
				end
				if(in == 3) begin
					state<=1084;
					out<=53;
				end
				if(in == 4) begin
					state<=4982;
					out<=54;
				end
			end
			3083: begin
				if(in == 0) begin
					state<=3084;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=6973;
					out<=57;
				end
				if(in == 3) begin
					state<=1085;
					out<=58;
				end
				if(in == 4) begin
					state<=4983;
					out<=59;
				end
			end
			3084: begin
				if(in == 0) begin
					state<=3085;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=6974;
					out<=62;
				end
				if(in == 3) begin
					state<=1086;
					out<=63;
				end
				if(in == 4) begin
					state<=4984;
					out<=64;
				end
			end
			3085: begin
				if(in == 0) begin
					state<=3086;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=6975;
					out<=67;
				end
				if(in == 3) begin
					state<=1087;
					out<=68;
				end
				if(in == 4) begin
					state<=4985;
					out<=69;
				end
			end
			3086: begin
				if(in == 0) begin
					state<=3087;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=6976;
					out<=72;
				end
				if(in == 3) begin
					state<=1088;
					out<=73;
				end
				if(in == 4) begin
					state<=4986;
					out<=74;
				end
			end
			3087: begin
				if(in == 0) begin
					state<=3088;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=6977;
					out<=77;
				end
				if(in == 3) begin
					state<=1089;
					out<=78;
				end
				if(in == 4) begin
					state<=4987;
					out<=79;
				end
			end
			3088: begin
				if(in == 0) begin
					state<=3089;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=6978;
					out<=82;
				end
				if(in == 3) begin
					state<=1090;
					out<=83;
				end
				if(in == 4) begin
					state<=4988;
					out<=84;
				end
			end
			3089: begin
				if(in == 0) begin
					state<=3090;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=6979;
					out<=87;
				end
				if(in == 3) begin
					state<=1091;
					out<=88;
				end
				if(in == 4) begin
					state<=4989;
					out<=89;
				end
			end
			3090: begin
				if(in == 0) begin
					state<=3091;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=6980;
					out<=92;
				end
				if(in == 3) begin
					state<=1092;
					out<=93;
				end
				if(in == 4) begin
					state<=4990;
					out<=94;
				end
			end
			3091: begin
				if(in == 0) begin
					state<=3092;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=6981;
					out<=97;
				end
				if(in == 3) begin
					state<=1093;
					out<=98;
				end
				if(in == 4) begin
					state<=4991;
					out<=99;
				end
			end
			3092: begin
				if(in == 0) begin
					state<=3093;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=6982;
					out<=102;
				end
				if(in == 3) begin
					state<=1094;
					out<=103;
				end
				if(in == 4) begin
					state<=4992;
					out<=104;
				end
			end
			3093: begin
				if(in == 0) begin
					state<=3094;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=6983;
					out<=107;
				end
				if(in == 3) begin
					state<=1095;
					out<=108;
				end
				if(in == 4) begin
					state<=4993;
					out<=109;
				end
			end
			3094: begin
				if(in == 0) begin
					state<=3095;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=6984;
					out<=112;
				end
				if(in == 3) begin
					state<=1096;
					out<=113;
				end
				if(in == 4) begin
					state<=4994;
					out<=114;
				end
			end
			3095: begin
				if(in == 0) begin
					state<=3096;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=6985;
					out<=117;
				end
				if(in == 3) begin
					state<=1097;
					out<=118;
				end
				if(in == 4) begin
					state<=4995;
					out<=119;
				end
			end
			3096: begin
				if(in == 0) begin
					state<=3097;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=6986;
					out<=122;
				end
				if(in == 3) begin
					state<=1098;
					out<=123;
				end
				if(in == 4) begin
					state<=4996;
					out<=124;
				end
			end
			3097: begin
				if(in == 0) begin
					state<=3098;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=6987;
					out<=127;
				end
				if(in == 3) begin
					state<=1099;
					out<=128;
				end
				if(in == 4) begin
					state<=4997;
					out<=129;
				end
			end
			3098: begin
				if(in == 0) begin
					state<=3099;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=6988;
					out<=132;
				end
				if(in == 3) begin
					state<=1100;
					out<=133;
				end
				if(in == 4) begin
					state<=4998;
					out<=134;
				end
			end
			3099: begin
				if(in == 0) begin
					state<=3100;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=6989;
					out<=137;
				end
				if(in == 3) begin
					state<=1101;
					out<=138;
				end
				if(in == 4) begin
					state<=4999;
					out<=139;
				end
			end
			3100: begin
				if(in == 0) begin
					state<=3101;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=6990;
					out<=142;
				end
				if(in == 3) begin
					state<=1102;
					out<=143;
				end
				if(in == 4) begin
					state<=5000;
					out<=144;
				end
			end
			3101: begin
				if(in == 0) begin
					state<=3102;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=6991;
					out<=147;
				end
				if(in == 3) begin
					state<=1103;
					out<=148;
				end
				if(in == 4) begin
					state<=5001;
					out<=149;
				end
			end
			3102: begin
				if(in == 0) begin
					state<=3103;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=6992;
					out<=152;
				end
				if(in == 3) begin
					state<=1104;
					out<=153;
				end
				if(in == 4) begin
					state<=5002;
					out<=154;
				end
			end
			3103: begin
				if(in == 0) begin
					state<=3104;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=6993;
					out<=157;
				end
				if(in == 3) begin
					state<=1105;
					out<=158;
				end
				if(in == 4) begin
					state<=5003;
					out<=159;
				end
			end
			3104: begin
				if(in == 0) begin
					state<=3105;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=6994;
					out<=162;
				end
				if(in == 3) begin
					state<=1106;
					out<=163;
				end
				if(in == 4) begin
					state<=5004;
					out<=164;
				end
			end
			3105: begin
				if(in == 0) begin
					state<=3106;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=6995;
					out<=167;
				end
				if(in == 3) begin
					state<=1107;
					out<=168;
				end
				if(in == 4) begin
					state<=5005;
					out<=169;
				end
			end
			3106: begin
				if(in == 0) begin
					state<=3107;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=6996;
					out<=172;
				end
				if(in == 3) begin
					state<=1108;
					out<=173;
				end
				if(in == 4) begin
					state<=5006;
					out<=174;
				end
			end
			3107: begin
				if(in == 0) begin
					state<=3108;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=6997;
					out<=177;
				end
				if(in == 3) begin
					state<=1109;
					out<=178;
				end
				if(in == 4) begin
					state<=5007;
					out<=179;
				end
			end
			3108: begin
				if(in == 0) begin
					state<=3109;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=6998;
					out<=182;
				end
				if(in == 3) begin
					state<=1110;
					out<=183;
				end
				if(in == 4) begin
					state<=5008;
					out<=184;
				end
			end
			3109: begin
				if(in == 0) begin
					state<=3110;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=6999;
					out<=187;
				end
				if(in == 3) begin
					state<=1111;
					out<=188;
				end
				if(in == 4) begin
					state<=5009;
					out<=189;
				end
			end
			3110: begin
				if(in == 0) begin
					state<=3111;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=7000;
					out<=192;
				end
				if(in == 3) begin
					state<=1112;
					out<=193;
				end
				if(in == 4) begin
					state<=5010;
					out<=194;
				end
			end
			3111: begin
				if(in == 0) begin
					state<=3112;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=7001;
					out<=197;
				end
				if(in == 3) begin
					state<=1113;
					out<=198;
				end
				if(in == 4) begin
					state<=5011;
					out<=199;
				end
			end
			3112: begin
				if(in == 0) begin
					state<=3113;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=7002;
					out<=202;
				end
				if(in == 3) begin
					state<=1114;
					out<=203;
				end
				if(in == 4) begin
					state<=5012;
					out<=204;
				end
			end
			3113: begin
				if(in == 0) begin
					state<=3114;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=7003;
					out<=207;
				end
				if(in == 3) begin
					state<=1115;
					out<=208;
				end
				if(in == 4) begin
					state<=5013;
					out<=209;
				end
			end
			3114: begin
				if(in == 0) begin
					state<=3115;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=7004;
					out<=212;
				end
				if(in == 3) begin
					state<=1116;
					out<=213;
				end
				if(in == 4) begin
					state<=5014;
					out<=214;
				end
			end
			3115: begin
				if(in == 0) begin
					state<=3116;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=7005;
					out<=217;
				end
				if(in == 3) begin
					state<=1117;
					out<=218;
				end
				if(in == 4) begin
					state<=5015;
					out<=219;
				end
			end
			3116: begin
				if(in == 0) begin
					state<=3117;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=7006;
					out<=222;
				end
				if(in == 3) begin
					state<=1118;
					out<=223;
				end
				if(in == 4) begin
					state<=5016;
					out<=224;
				end
			end
			3117: begin
				if(in == 0) begin
					state<=3118;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=7007;
					out<=227;
				end
				if(in == 3) begin
					state<=1119;
					out<=228;
				end
				if(in == 4) begin
					state<=5017;
					out<=229;
				end
			end
			3118: begin
				if(in == 0) begin
					state<=3119;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=7008;
					out<=232;
				end
				if(in == 3) begin
					state<=1120;
					out<=233;
				end
				if(in == 4) begin
					state<=5018;
					out<=234;
				end
			end
			3119: begin
				if(in == 0) begin
					state<=3120;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=7009;
					out<=237;
				end
				if(in == 3) begin
					state<=1121;
					out<=238;
				end
				if(in == 4) begin
					state<=5019;
					out<=239;
				end
			end
			3120: begin
				if(in == 0) begin
					state<=3121;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=7010;
					out<=242;
				end
				if(in == 3) begin
					state<=1122;
					out<=243;
				end
				if(in == 4) begin
					state<=5020;
					out<=244;
				end
			end
			3121: begin
				if(in == 0) begin
					state<=3122;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=7011;
					out<=247;
				end
				if(in == 3) begin
					state<=1123;
					out<=248;
				end
				if(in == 4) begin
					state<=5021;
					out<=249;
				end
			end
			3122: begin
				if(in == 0) begin
					state<=3123;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=7012;
					out<=252;
				end
				if(in == 3) begin
					state<=1124;
					out<=253;
				end
				if(in == 4) begin
					state<=5022;
					out<=254;
				end
			end
			3123: begin
				if(in == 0) begin
					state<=3124;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=7013;
					out<=1;
				end
				if(in == 3) begin
					state<=1125;
					out<=2;
				end
				if(in == 4) begin
					state<=5023;
					out<=3;
				end
			end
			3124: begin
				if(in == 0) begin
					state<=3125;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=7014;
					out<=6;
				end
				if(in == 3) begin
					state<=1126;
					out<=7;
				end
				if(in == 4) begin
					state<=5024;
					out<=8;
				end
			end
			3125: begin
				if(in == 0) begin
					state<=3126;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=7015;
					out<=11;
				end
				if(in == 3) begin
					state<=1127;
					out<=12;
				end
				if(in == 4) begin
					state<=5025;
					out<=13;
				end
			end
			3126: begin
				if(in == 0) begin
					state<=3127;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=7016;
					out<=16;
				end
				if(in == 3) begin
					state<=1128;
					out<=17;
				end
				if(in == 4) begin
					state<=5026;
					out<=18;
				end
			end
			3127: begin
				if(in == 0) begin
					state<=3128;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=7017;
					out<=21;
				end
				if(in == 3) begin
					state<=1129;
					out<=22;
				end
				if(in == 4) begin
					state<=5027;
					out<=23;
				end
			end
			3128: begin
				if(in == 0) begin
					state<=3129;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=7018;
					out<=26;
				end
				if(in == 3) begin
					state<=1130;
					out<=27;
				end
				if(in == 4) begin
					state<=5028;
					out<=28;
				end
			end
			3129: begin
				if(in == 0) begin
					state<=3130;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=7019;
					out<=31;
				end
				if(in == 3) begin
					state<=1131;
					out<=32;
				end
				if(in == 4) begin
					state<=5029;
					out<=33;
				end
			end
			3130: begin
				if(in == 0) begin
					state<=3131;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=7020;
					out<=36;
				end
				if(in == 3) begin
					state<=1132;
					out<=37;
				end
				if(in == 4) begin
					state<=5030;
					out<=38;
				end
			end
			3131: begin
				if(in == 0) begin
					state<=3132;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=7021;
					out<=41;
				end
				if(in == 3) begin
					state<=1133;
					out<=42;
				end
				if(in == 4) begin
					state<=5031;
					out<=43;
				end
			end
			3132: begin
				if(in == 0) begin
					state<=3133;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=7022;
					out<=46;
				end
				if(in == 3) begin
					state<=1134;
					out<=47;
				end
				if(in == 4) begin
					state<=5032;
					out<=48;
				end
			end
			3133: begin
				if(in == 0) begin
					state<=3134;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=7023;
					out<=51;
				end
				if(in == 3) begin
					state<=1135;
					out<=52;
				end
				if(in == 4) begin
					state<=5033;
					out<=53;
				end
			end
			3134: begin
				if(in == 0) begin
					state<=3135;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=7024;
					out<=56;
				end
				if(in == 3) begin
					state<=1136;
					out<=57;
				end
				if(in == 4) begin
					state<=5034;
					out<=58;
				end
			end
			3135: begin
				if(in == 0) begin
					state<=3136;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=7025;
					out<=61;
				end
				if(in == 3) begin
					state<=1137;
					out<=62;
				end
				if(in == 4) begin
					state<=5035;
					out<=63;
				end
			end
			3136: begin
				if(in == 0) begin
					state<=3137;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=7026;
					out<=66;
				end
				if(in == 3) begin
					state<=1138;
					out<=67;
				end
				if(in == 4) begin
					state<=5036;
					out<=68;
				end
			end
			3137: begin
				if(in == 0) begin
					state<=3138;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=7027;
					out<=71;
				end
				if(in == 3) begin
					state<=1139;
					out<=72;
				end
				if(in == 4) begin
					state<=5037;
					out<=73;
				end
			end
			3138: begin
				if(in == 0) begin
					state<=3139;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=7028;
					out<=76;
				end
				if(in == 3) begin
					state<=1140;
					out<=77;
				end
				if(in == 4) begin
					state<=5038;
					out<=78;
				end
			end
			3139: begin
				if(in == 0) begin
					state<=3140;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=7029;
					out<=81;
				end
				if(in == 3) begin
					state<=1141;
					out<=82;
				end
				if(in == 4) begin
					state<=5039;
					out<=83;
				end
			end
			3140: begin
				if(in == 0) begin
					state<=3141;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=7030;
					out<=86;
				end
				if(in == 3) begin
					state<=1142;
					out<=87;
				end
				if(in == 4) begin
					state<=5040;
					out<=88;
				end
			end
			3141: begin
				if(in == 0) begin
					state<=3142;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=7031;
					out<=91;
				end
				if(in == 3) begin
					state<=1143;
					out<=92;
				end
				if(in == 4) begin
					state<=5041;
					out<=93;
				end
			end
			3142: begin
				if(in == 0) begin
					state<=3143;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=7032;
					out<=96;
				end
				if(in == 3) begin
					state<=1144;
					out<=97;
				end
				if(in == 4) begin
					state<=5042;
					out<=98;
				end
			end
			3143: begin
				if(in == 0) begin
					state<=3144;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=7033;
					out<=101;
				end
				if(in == 3) begin
					state<=1145;
					out<=102;
				end
				if(in == 4) begin
					state<=5043;
					out<=103;
				end
			end
			3144: begin
				if(in == 0) begin
					state<=3145;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=7034;
					out<=106;
				end
				if(in == 3) begin
					state<=1146;
					out<=107;
				end
				if(in == 4) begin
					state<=5044;
					out<=108;
				end
			end
			3145: begin
				if(in == 0) begin
					state<=3146;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=7035;
					out<=111;
				end
				if(in == 3) begin
					state<=1147;
					out<=112;
				end
				if(in == 4) begin
					state<=5045;
					out<=113;
				end
			end
			3146: begin
				if(in == 0) begin
					state<=3147;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=7036;
					out<=116;
				end
				if(in == 3) begin
					state<=1148;
					out<=117;
				end
				if(in == 4) begin
					state<=5046;
					out<=118;
				end
			end
			3147: begin
				if(in == 0) begin
					state<=3148;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=7037;
					out<=121;
				end
				if(in == 3) begin
					state<=1149;
					out<=122;
				end
				if(in == 4) begin
					state<=5047;
					out<=123;
				end
			end
			3148: begin
				if(in == 0) begin
					state<=3149;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=7038;
					out<=126;
				end
				if(in == 3) begin
					state<=1150;
					out<=127;
				end
				if(in == 4) begin
					state<=5048;
					out<=128;
				end
			end
			3149: begin
				if(in == 0) begin
					state<=3150;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=7039;
					out<=131;
				end
				if(in == 3) begin
					state<=1151;
					out<=132;
				end
				if(in == 4) begin
					state<=5049;
					out<=133;
				end
			end
			3150: begin
				if(in == 0) begin
					state<=3151;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=7040;
					out<=136;
				end
				if(in == 3) begin
					state<=1152;
					out<=137;
				end
				if(in == 4) begin
					state<=5050;
					out<=138;
				end
			end
			3151: begin
				if(in == 0) begin
					state<=3152;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=7041;
					out<=141;
				end
				if(in == 3) begin
					state<=1153;
					out<=142;
				end
				if(in == 4) begin
					state<=5051;
					out<=143;
				end
			end
			3152: begin
				if(in == 0) begin
					state<=3153;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=7042;
					out<=146;
				end
				if(in == 3) begin
					state<=1154;
					out<=147;
				end
				if(in == 4) begin
					state<=5052;
					out<=148;
				end
			end
			3153: begin
				if(in == 0) begin
					state<=3154;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=7043;
					out<=151;
				end
				if(in == 3) begin
					state<=1155;
					out<=152;
				end
				if(in == 4) begin
					state<=5053;
					out<=153;
				end
			end
			3154: begin
				if(in == 0) begin
					state<=3155;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=7044;
					out<=156;
				end
				if(in == 3) begin
					state<=1156;
					out<=157;
				end
				if(in == 4) begin
					state<=5054;
					out<=158;
				end
			end
			3155: begin
				if(in == 0) begin
					state<=3156;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=7045;
					out<=161;
				end
				if(in == 3) begin
					state<=1157;
					out<=162;
				end
				if(in == 4) begin
					state<=5055;
					out<=163;
				end
			end
			3156: begin
				if(in == 0) begin
					state<=3157;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=7046;
					out<=166;
				end
				if(in == 3) begin
					state<=1158;
					out<=167;
				end
				if(in == 4) begin
					state<=5056;
					out<=168;
				end
			end
			3157: begin
				if(in == 0) begin
					state<=3158;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=7047;
					out<=171;
				end
				if(in == 3) begin
					state<=1159;
					out<=172;
				end
				if(in == 4) begin
					state<=5057;
					out<=173;
				end
			end
			3158: begin
				if(in == 0) begin
					state<=3159;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=7048;
					out<=176;
				end
				if(in == 3) begin
					state<=1160;
					out<=177;
				end
				if(in == 4) begin
					state<=5058;
					out<=178;
				end
			end
			3159: begin
				if(in == 0) begin
					state<=3160;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=7049;
					out<=181;
				end
				if(in == 3) begin
					state<=1161;
					out<=182;
				end
				if(in == 4) begin
					state<=5059;
					out<=183;
				end
			end
			3160: begin
				if(in == 0) begin
					state<=3161;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=7050;
					out<=186;
				end
				if(in == 3) begin
					state<=1162;
					out<=187;
				end
				if(in == 4) begin
					state<=5060;
					out<=188;
				end
			end
			3161: begin
				if(in == 0) begin
					state<=3162;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=7051;
					out<=191;
				end
				if(in == 3) begin
					state<=1163;
					out<=192;
				end
				if(in == 4) begin
					state<=5061;
					out<=193;
				end
			end
			3162: begin
				if(in == 0) begin
					state<=3163;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=7052;
					out<=196;
				end
				if(in == 3) begin
					state<=1164;
					out<=197;
				end
				if(in == 4) begin
					state<=5062;
					out<=198;
				end
			end
			3163: begin
				if(in == 0) begin
					state<=3164;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=7053;
					out<=201;
				end
				if(in == 3) begin
					state<=1165;
					out<=202;
				end
				if(in == 4) begin
					state<=5063;
					out<=203;
				end
			end
			3164: begin
				if(in == 0) begin
					state<=3165;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=7054;
					out<=206;
				end
				if(in == 3) begin
					state<=1166;
					out<=207;
				end
				if(in == 4) begin
					state<=5064;
					out<=208;
				end
			end
			3165: begin
				if(in == 0) begin
					state<=3166;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=7055;
					out<=211;
				end
				if(in == 3) begin
					state<=1167;
					out<=212;
				end
				if(in == 4) begin
					state<=5065;
					out<=213;
				end
			end
			3166: begin
				if(in == 0) begin
					state<=3167;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=7056;
					out<=216;
				end
				if(in == 3) begin
					state<=1168;
					out<=217;
				end
				if(in == 4) begin
					state<=5066;
					out<=218;
				end
			end
			3167: begin
				if(in == 0) begin
					state<=3168;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=7057;
					out<=221;
				end
				if(in == 3) begin
					state<=1169;
					out<=222;
				end
				if(in == 4) begin
					state<=5067;
					out<=223;
				end
			end
			3168: begin
				if(in == 0) begin
					state<=3169;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=7058;
					out<=226;
				end
				if(in == 3) begin
					state<=1170;
					out<=227;
				end
				if(in == 4) begin
					state<=5068;
					out<=228;
				end
			end
			3169: begin
				if(in == 0) begin
					state<=3170;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=7059;
					out<=231;
				end
				if(in == 3) begin
					state<=1171;
					out<=232;
				end
				if(in == 4) begin
					state<=5069;
					out<=233;
				end
			end
			3170: begin
				if(in == 0) begin
					state<=3171;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=7060;
					out<=236;
				end
				if(in == 3) begin
					state<=1172;
					out<=237;
				end
				if(in == 4) begin
					state<=5070;
					out<=238;
				end
			end
			3171: begin
				if(in == 0) begin
					state<=3172;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=7061;
					out<=241;
				end
				if(in == 3) begin
					state<=1173;
					out<=242;
				end
				if(in == 4) begin
					state<=5071;
					out<=243;
				end
			end
			3172: begin
				if(in == 0) begin
					state<=3173;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=7062;
					out<=246;
				end
				if(in == 3) begin
					state<=1174;
					out<=247;
				end
				if(in == 4) begin
					state<=5072;
					out<=248;
				end
			end
			3173: begin
				if(in == 0) begin
					state<=3174;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=7063;
					out<=251;
				end
				if(in == 3) begin
					state<=1175;
					out<=252;
				end
				if(in == 4) begin
					state<=5073;
					out<=253;
				end
			end
			3174: begin
				if(in == 0) begin
					state<=3175;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=7064;
					out<=0;
				end
				if(in == 3) begin
					state<=1176;
					out<=1;
				end
				if(in == 4) begin
					state<=5074;
					out<=2;
				end
			end
			3175: begin
				if(in == 0) begin
					state<=3176;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=7065;
					out<=5;
				end
				if(in == 3) begin
					state<=1177;
					out<=6;
				end
				if(in == 4) begin
					state<=5075;
					out<=7;
				end
			end
			3176: begin
				if(in == 0) begin
					state<=3177;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=7066;
					out<=10;
				end
				if(in == 3) begin
					state<=1178;
					out<=11;
				end
				if(in == 4) begin
					state<=5076;
					out<=12;
				end
			end
			3177: begin
				if(in == 0) begin
					state<=3178;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=7067;
					out<=15;
				end
				if(in == 3) begin
					state<=1179;
					out<=16;
				end
				if(in == 4) begin
					state<=5077;
					out<=17;
				end
			end
			3178: begin
				if(in == 0) begin
					state<=3179;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=7068;
					out<=20;
				end
				if(in == 3) begin
					state<=1180;
					out<=21;
				end
				if(in == 4) begin
					state<=5078;
					out<=22;
				end
			end
			3179: begin
				if(in == 0) begin
					state<=3180;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=7069;
					out<=25;
				end
				if(in == 3) begin
					state<=1181;
					out<=26;
				end
				if(in == 4) begin
					state<=5079;
					out<=27;
				end
			end
			3180: begin
				if(in == 0) begin
					state<=3181;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=7070;
					out<=30;
				end
				if(in == 3) begin
					state<=1182;
					out<=31;
				end
				if(in == 4) begin
					state<=5080;
					out<=32;
				end
			end
			3181: begin
				if(in == 0) begin
					state<=3182;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=7071;
					out<=35;
				end
				if(in == 3) begin
					state<=1183;
					out<=36;
				end
				if(in == 4) begin
					state<=5081;
					out<=37;
				end
			end
			3182: begin
				if(in == 0) begin
					state<=3183;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=7072;
					out<=40;
				end
				if(in == 3) begin
					state<=1184;
					out<=41;
				end
				if(in == 4) begin
					state<=5082;
					out<=42;
				end
			end
			3183: begin
				if(in == 0) begin
					state<=3184;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=7073;
					out<=45;
				end
				if(in == 3) begin
					state<=1185;
					out<=46;
				end
				if(in == 4) begin
					state<=5083;
					out<=47;
				end
			end
			3184: begin
				if(in == 0) begin
					state<=3185;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=7074;
					out<=50;
				end
				if(in == 3) begin
					state<=1186;
					out<=51;
				end
				if(in == 4) begin
					state<=5084;
					out<=52;
				end
			end
			3185: begin
				if(in == 0) begin
					state<=3186;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=7075;
					out<=55;
				end
				if(in == 3) begin
					state<=1187;
					out<=56;
				end
				if(in == 4) begin
					state<=5085;
					out<=57;
				end
			end
			3186: begin
				if(in == 0) begin
					state<=3187;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=7076;
					out<=60;
				end
				if(in == 3) begin
					state<=1188;
					out<=61;
				end
				if(in == 4) begin
					state<=5086;
					out<=62;
				end
			end
			3187: begin
				if(in == 0) begin
					state<=3188;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=7077;
					out<=65;
				end
				if(in == 3) begin
					state<=1189;
					out<=66;
				end
				if(in == 4) begin
					state<=5087;
					out<=67;
				end
			end
			3188: begin
				if(in == 0) begin
					state<=3189;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=7078;
					out<=70;
				end
				if(in == 3) begin
					state<=1190;
					out<=71;
				end
				if(in == 4) begin
					state<=5088;
					out<=72;
				end
			end
			3189: begin
				if(in == 0) begin
					state<=3190;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=7079;
					out<=75;
				end
				if(in == 3) begin
					state<=1191;
					out<=76;
				end
				if(in == 4) begin
					state<=5089;
					out<=77;
				end
			end
			3190: begin
				if(in == 0) begin
					state<=3191;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=7080;
					out<=80;
				end
				if(in == 3) begin
					state<=1192;
					out<=81;
				end
				if(in == 4) begin
					state<=5090;
					out<=82;
				end
			end
			3191: begin
				if(in == 0) begin
					state<=3192;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=7081;
					out<=85;
				end
				if(in == 3) begin
					state<=1193;
					out<=86;
				end
				if(in == 4) begin
					state<=5091;
					out<=87;
				end
			end
			3192: begin
				if(in == 0) begin
					state<=3193;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=7082;
					out<=90;
				end
				if(in == 3) begin
					state<=1194;
					out<=91;
				end
				if(in == 4) begin
					state<=5092;
					out<=92;
				end
			end
			3193: begin
				if(in == 0) begin
					state<=3194;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=7083;
					out<=95;
				end
				if(in == 3) begin
					state<=1195;
					out<=96;
				end
				if(in == 4) begin
					state<=5093;
					out<=97;
				end
			end
			3194: begin
				if(in == 0) begin
					state<=3195;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=7084;
					out<=100;
				end
				if(in == 3) begin
					state<=1196;
					out<=101;
				end
				if(in == 4) begin
					state<=5094;
					out<=102;
				end
			end
			3195: begin
				if(in == 0) begin
					state<=3196;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=7085;
					out<=105;
				end
				if(in == 3) begin
					state<=1197;
					out<=106;
				end
				if(in == 4) begin
					state<=5095;
					out<=107;
				end
			end
			3196: begin
				if(in == 0) begin
					state<=3197;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=7086;
					out<=110;
				end
				if(in == 3) begin
					state<=1198;
					out<=111;
				end
				if(in == 4) begin
					state<=5096;
					out<=112;
				end
			end
			3197: begin
				if(in == 0) begin
					state<=3198;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=7087;
					out<=115;
				end
				if(in == 3) begin
					state<=1199;
					out<=116;
				end
				if(in == 4) begin
					state<=5097;
					out<=117;
				end
			end
			3198: begin
				if(in == 0) begin
					state<=3199;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=7088;
					out<=120;
				end
				if(in == 3) begin
					state<=1200;
					out<=121;
				end
				if(in == 4) begin
					state<=5098;
					out<=122;
				end
			end
			3199: begin
				if(in == 0) begin
					state<=3200;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=7089;
					out<=125;
				end
				if(in == 3) begin
					state<=1201;
					out<=126;
				end
				if(in == 4) begin
					state<=5099;
					out<=127;
				end
			end
			3200: begin
				if(in == 0) begin
					state<=3201;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=7090;
					out<=130;
				end
				if(in == 3) begin
					state<=1202;
					out<=131;
				end
				if(in == 4) begin
					state<=5100;
					out<=132;
				end
			end
			3201: begin
				if(in == 0) begin
					state<=3202;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=7091;
					out<=135;
				end
				if(in == 3) begin
					state<=1203;
					out<=136;
				end
				if(in == 4) begin
					state<=5101;
					out<=137;
				end
			end
			3202: begin
				if(in == 0) begin
					state<=3203;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=7092;
					out<=140;
				end
				if(in == 3) begin
					state<=1204;
					out<=141;
				end
				if(in == 4) begin
					state<=5102;
					out<=142;
				end
			end
			3203: begin
				if(in == 0) begin
					state<=3204;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=7093;
					out<=145;
				end
				if(in == 3) begin
					state<=1205;
					out<=146;
				end
				if(in == 4) begin
					state<=5103;
					out<=147;
				end
			end
			3204: begin
				if(in == 0) begin
					state<=3205;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=7094;
					out<=150;
				end
				if(in == 3) begin
					state<=1206;
					out<=151;
				end
				if(in == 4) begin
					state<=5104;
					out<=152;
				end
			end
			3205: begin
				if(in == 0) begin
					state<=3206;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=7095;
					out<=155;
				end
				if(in == 3) begin
					state<=1207;
					out<=156;
				end
				if(in == 4) begin
					state<=5105;
					out<=157;
				end
			end
			3206: begin
				if(in == 0) begin
					state<=3207;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=7096;
					out<=160;
				end
				if(in == 3) begin
					state<=1208;
					out<=161;
				end
				if(in == 4) begin
					state<=5106;
					out<=162;
				end
			end
			3207: begin
				if(in == 0) begin
					state<=3208;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=7097;
					out<=165;
				end
				if(in == 3) begin
					state<=1209;
					out<=166;
				end
				if(in == 4) begin
					state<=5107;
					out<=167;
				end
			end
			3208: begin
				if(in == 0) begin
					state<=3209;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=7098;
					out<=170;
				end
				if(in == 3) begin
					state<=1210;
					out<=171;
				end
				if(in == 4) begin
					state<=5108;
					out<=172;
				end
			end
			3209: begin
				if(in == 0) begin
					state<=3210;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=7099;
					out<=175;
				end
				if(in == 3) begin
					state<=1211;
					out<=176;
				end
				if(in == 4) begin
					state<=5109;
					out<=177;
				end
			end
			3210: begin
				if(in == 0) begin
					state<=3211;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=7100;
					out<=180;
				end
				if(in == 3) begin
					state<=1212;
					out<=181;
				end
				if(in == 4) begin
					state<=5110;
					out<=182;
				end
			end
			3211: begin
				if(in == 0) begin
					state<=3212;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=7101;
					out<=185;
				end
				if(in == 3) begin
					state<=1213;
					out<=186;
				end
				if(in == 4) begin
					state<=5111;
					out<=187;
				end
			end
			3212: begin
				if(in == 0) begin
					state<=3213;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=7102;
					out<=190;
				end
				if(in == 3) begin
					state<=1214;
					out<=191;
				end
				if(in == 4) begin
					state<=5112;
					out<=192;
				end
			end
			3213: begin
				if(in == 0) begin
					state<=3214;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=7103;
					out<=195;
				end
				if(in == 3) begin
					state<=1215;
					out<=196;
				end
				if(in == 4) begin
					state<=5113;
					out<=197;
				end
			end
			3214: begin
				if(in == 0) begin
					state<=3215;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=7104;
					out<=200;
				end
				if(in == 3) begin
					state<=1216;
					out<=201;
				end
				if(in == 4) begin
					state<=5114;
					out<=202;
				end
			end
			3215: begin
				if(in == 0) begin
					state<=3216;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=7105;
					out<=205;
				end
				if(in == 3) begin
					state<=1217;
					out<=206;
				end
				if(in == 4) begin
					state<=5115;
					out<=207;
				end
			end
			3216: begin
				if(in == 0) begin
					state<=3217;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=7106;
					out<=210;
				end
				if(in == 3) begin
					state<=1218;
					out<=211;
				end
				if(in == 4) begin
					state<=5116;
					out<=212;
				end
			end
			3217: begin
				if(in == 0) begin
					state<=3218;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=7107;
					out<=215;
				end
				if(in == 3) begin
					state<=1219;
					out<=216;
				end
				if(in == 4) begin
					state<=5117;
					out<=217;
				end
			end
			3218: begin
				if(in == 0) begin
					state<=3219;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=7108;
					out<=220;
				end
				if(in == 3) begin
					state<=1220;
					out<=221;
				end
				if(in == 4) begin
					state<=5118;
					out<=222;
				end
			end
			3219: begin
				if(in == 0) begin
					state<=3220;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=7109;
					out<=225;
				end
				if(in == 3) begin
					state<=1221;
					out<=226;
				end
				if(in == 4) begin
					state<=5119;
					out<=227;
				end
			end
			3220: begin
				if(in == 0) begin
					state<=3221;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=7110;
					out<=230;
				end
				if(in == 3) begin
					state<=1222;
					out<=231;
				end
				if(in == 4) begin
					state<=5120;
					out<=232;
				end
			end
			3221: begin
				if(in == 0) begin
					state<=3222;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=7111;
					out<=235;
				end
				if(in == 3) begin
					state<=1223;
					out<=236;
				end
				if(in == 4) begin
					state<=5121;
					out<=237;
				end
			end
			3222: begin
				if(in == 0) begin
					state<=3223;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=7112;
					out<=240;
				end
				if(in == 3) begin
					state<=1224;
					out<=241;
				end
				if(in == 4) begin
					state<=5122;
					out<=242;
				end
			end
			3223: begin
				if(in == 0) begin
					state<=3224;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=7113;
					out<=245;
				end
				if(in == 3) begin
					state<=1225;
					out<=246;
				end
				if(in == 4) begin
					state<=5123;
					out<=247;
				end
			end
			3224: begin
				if(in == 0) begin
					state<=3225;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=7114;
					out<=250;
				end
				if(in == 3) begin
					state<=1226;
					out<=251;
				end
				if(in == 4) begin
					state<=5124;
					out<=252;
				end
			end
			3225: begin
				if(in == 0) begin
					state<=3226;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=7115;
					out<=255;
				end
				if(in == 3) begin
					state<=1227;
					out<=0;
				end
				if(in == 4) begin
					state<=5125;
					out<=1;
				end
			end
			3226: begin
				if(in == 0) begin
					state<=3227;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=7116;
					out<=4;
				end
				if(in == 3) begin
					state<=1228;
					out<=5;
				end
				if(in == 4) begin
					state<=5126;
					out<=6;
				end
			end
			3227: begin
				if(in == 0) begin
					state<=3228;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=7117;
					out<=9;
				end
				if(in == 3) begin
					state<=1229;
					out<=10;
				end
				if(in == 4) begin
					state<=5127;
					out<=11;
				end
			end
			3228: begin
				if(in == 0) begin
					state<=3229;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=7118;
					out<=14;
				end
				if(in == 3) begin
					state<=1230;
					out<=15;
				end
				if(in == 4) begin
					state<=5128;
					out<=16;
				end
			end
			3229: begin
				if(in == 0) begin
					state<=2689;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=6578;
					out<=19;
				end
				if(in == 3) begin
					state<=691;
					out<=20;
				end
				if(in == 4) begin
					state<=4589;
					out<=21;
				end
			end
			3230: begin
				if(in == 0) begin
					state<=3231;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=7120;
					out<=24;
				end
				if(in == 3) begin
					state<=1578;
					out<=25;
				end
				if(in == 4) begin
					state<=5467;
					out<=26;
				end
			end
			3231: begin
				if(in == 0) begin
					state<=3232;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=7121;
					out<=29;
				end
				if(in == 3) begin
					state<=1579;
					out<=30;
				end
				if(in == 4) begin
					state<=5468;
					out<=31;
				end
			end
			3232: begin
				if(in == 0) begin
					state<=3233;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=7122;
					out<=34;
				end
				if(in == 3) begin
					state<=1580;
					out<=35;
				end
				if(in == 4) begin
					state<=5469;
					out<=36;
				end
			end
			3233: begin
				if(in == 0) begin
					state<=3234;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=7123;
					out<=39;
				end
				if(in == 3) begin
					state<=1581;
					out<=40;
				end
				if(in == 4) begin
					state<=5470;
					out<=41;
				end
			end
			3234: begin
				if(in == 0) begin
					state<=3235;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=7124;
					out<=44;
				end
				if(in == 3) begin
					state<=1582;
					out<=45;
				end
				if(in == 4) begin
					state<=5471;
					out<=46;
				end
			end
			3235: begin
				if(in == 0) begin
					state<=3236;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=7125;
					out<=49;
				end
				if(in == 3) begin
					state<=1583;
					out<=50;
				end
				if(in == 4) begin
					state<=5472;
					out<=51;
				end
			end
			3236: begin
				if(in == 0) begin
					state<=3237;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=7126;
					out<=54;
				end
				if(in == 3) begin
					state<=1584;
					out<=55;
				end
				if(in == 4) begin
					state<=5473;
					out<=56;
				end
			end
			3237: begin
				if(in == 0) begin
					state<=3238;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=7127;
					out<=59;
				end
				if(in == 3) begin
					state<=1585;
					out<=60;
				end
				if(in == 4) begin
					state<=5474;
					out<=61;
				end
			end
			3238: begin
				if(in == 0) begin
					state<=3239;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=7128;
					out<=64;
				end
				if(in == 3) begin
					state<=1586;
					out<=65;
				end
				if(in == 4) begin
					state<=5475;
					out<=66;
				end
			end
			3239: begin
				if(in == 0) begin
					state<=3240;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=7129;
					out<=69;
				end
				if(in == 3) begin
					state<=1587;
					out<=70;
				end
				if(in == 4) begin
					state<=5476;
					out<=71;
				end
			end
			3240: begin
				if(in == 0) begin
					state<=3241;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=7130;
					out<=74;
				end
				if(in == 3) begin
					state<=1588;
					out<=75;
				end
				if(in == 4) begin
					state<=5477;
					out<=76;
				end
			end
			3241: begin
				if(in == 0) begin
					state<=3242;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=7131;
					out<=79;
				end
				if(in == 3) begin
					state<=1589;
					out<=80;
				end
				if(in == 4) begin
					state<=5478;
					out<=81;
				end
			end
			3242: begin
				if(in == 0) begin
					state<=3243;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=7132;
					out<=84;
				end
				if(in == 3) begin
					state<=1590;
					out<=85;
				end
				if(in == 4) begin
					state<=5479;
					out<=86;
				end
			end
			3243: begin
				if(in == 0) begin
					state<=3244;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=7133;
					out<=89;
				end
				if(in == 3) begin
					state<=1591;
					out<=90;
				end
				if(in == 4) begin
					state<=5480;
					out<=91;
				end
			end
			3244: begin
				if(in == 0) begin
					state<=3245;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=7134;
					out<=94;
				end
				if(in == 3) begin
					state<=1592;
					out<=95;
				end
				if(in == 4) begin
					state<=5481;
					out<=96;
				end
			end
			3245: begin
				if(in == 0) begin
					state<=3246;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=7135;
					out<=99;
				end
				if(in == 3) begin
					state<=1593;
					out<=100;
				end
				if(in == 4) begin
					state<=5482;
					out<=101;
				end
			end
			3246: begin
				if(in == 0) begin
					state<=3247;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=7136;
					out<=104;
				end
				if(in == 3) begin
					state<=1594;
					out<=105;
				end
				if(in == 4) begin
					state<=5483;
					out<=106;
				end
			end
			3247: begin
				if(in == 0) begin
					state<=3248;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=7137;
					out<=109;
				end
				if(in == 3) begin
					state<=1595;
					out<=110;
				end
				if(in == 4) begin
					state<=5484;
					out<=111;
				end
			end
			3248: begin
				if(in == 0) begin
					state<=3249;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=7138;
					out<=114;
				end
				if(in == 3) begin
					state<=1596;
					out<=115;
				end
				if(in == 4) begin
					state<=5485;
					out<=116;
				end
			end
			3249: begin
				if(in == 0) begin
					state<=3250;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=7139;
					out<=119;
				end
				if(in == 3) begin
					state<=1597;
					out<=120;
				end
				if(in == 4) begin
					state<=5486;
					out<=121;
				end
			end
			3250: begin
				if(in == 0) begin
					state<=3251;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=7140;
					out<=124;
				end
				if(in == 3) begin
					state<=1598;
					out<=125;
				end
				if(in == 4) begin
					state<=5487;
					out<=126;
				end
			end
			3251: begin
				if(in == 0) begin
					state<=3252;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=7141;
					out<=129;
				end
				if(in == 3) begin
					state<=1599;
					out<=130;
				end
				if(in == 4) begin
					state<=5488;
					out<=131;
				end
			end
			3252: begin
				if(in == 0) begin
					state<=3253;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=7142;
					out<=134;
				end
				if(in == 3) begin
					state<=1600;
					out<=135;
				end
				if(in == 4) begin
					state<=5489;
					out<=136;
				end
			end
			3253: begin
				if(in == 0) begin
					state<=3254;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=7143;
					out<=139;
				end
				if(in == 3) begin
					state<=1601;
					out<=140;
				end
				if(in == 4) begin
					state<=5490;
					out<=141;
				end
			end
			3254: begin
				if(in == 0) begin
					state<=3255;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=7144;
					out<=144;
				end
				if(in == 3) begin
					state<=1602;
					out<=145;
				end
				if(in == 4) begin
					state<=5491;
					out<=146;
				end
			end
			3255: begin
				if(in == 0) begin
					state<=3256;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=7145;
					out<=149;
				end
				if(in == 3) begin
					state<=1603;
					out<=150;
				end
				if(in == 4) begin
					state<=5492;
					out<=151;
				end
			end
			3256: begin
				if(in == 0) begin
					state<=3257;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=7146;
					out<=154;
				end
				if(in == 3) begin
					state<=1604;
					out<=155;
				end
				if(in == 4) begin
					state<=5493;
					out<=156;
				end
			end
			3257: begin
				if(in == 0) begin
					state<=3258;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=7147;
					out<=159;
				end
				if(in == 3) begin
					state<=1605;
					out<=160;
				end
				if(in == 4) begin
					state<=5494;
					out<=161;
				end
			end
			3258: begin
				if(in == 0) begin
					state<=3259;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=7148;
					out<=164;
				end
				if(in == 3) begin
					state<=1606;
					out<=165;
				end
				if(in == 4) begin
					state<=5495;
					out<=166;
				end
			end
			3259: begin
				if(in == 0) begin
					state<=3260;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=7149;
					out<=169;
				end
				if(in == 3) begin
					state<=1607;
					out<=170;
				end
				if(in == 4) begin
					state<=5496;
					out<=171;
				end
			end
			3260: begin
				if(in == 0) begin
					state<=2670;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=6559;
					out<=174;
				end
				if(in == 3) begin
					state<=672;
					out<=175;
				end
				if(in == 4) begin
					state<=4570;
					out<=176;
				end
			end
			3261: begin
				if(in == 0) begin
					state<=3262;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=7151;
					out<=179;
				end
				if(in == 3) begin
					state<=1330;
					out<=180;
				end
				if(in == 4) begin
					state<=5219;
					out<=181;
				end
			end
			3262: begin
				if(in == 0) begin
					state<=3263;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=7152;
					out<=184;
				end
				if(in == 3) begin
					state<=1331;
					out<=185;
				end
				if(in == 4) begin
					state<=5220;
					out<=186;
				end
			end
			3263: begin
				if(in == 0) begin
					state<=3264;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=7153;
					out<=189;
				end
				if(in == 3) begin
					state<=1332;
					out<=190;
				end
				if(in == 4) begin
					state<=5221;
					out<=191;
				end
			end
			3264: begin
				if(in == 0) begin
					state<=3265;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=7154;
					out<=194;
				end
				if(in == 3) begin
					state<=1333;
					out<=195;
				end
				if(in == 4) begin
					state<=5222;
					out<=196;
				end
			end
			3265: begin
				if(in == 0) begin
					state<=3266;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=7155;
					out<=199;
				end
				if(in == 3) begin
					state<=1334;
					out<=200;
				end
				if(in == 4) begin
					state<=5223;
					out<=201;
				end
			end
			3266: begin
				if(in == 0) begin
					state<=3267;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=7156;
					out<=204;
				end
				if(in == 3) begin
					state<=1335;
					out<=205;
				end
				if(in == 4) begin
					state<=5224;
					out<=206;
				end
			end
			3267: begin
				if(in == 0) begin
					state<=3268;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=7157;
					out<=209;
				end
				if(in == 3) begin
					state<=1336;
					out<=210;
				end
				if(in == 4) begin
					state<=5225;
					out<=211;
				end
			end
			3268: begin
				if(in == 0) begin
					state<=3269;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=7158;
					out<=214;
				end
				if(in == 3) begin
					state<=1337;
					out<=215;
				end
				if(in == 4) begin
					state<=5226;
					out<=216;
				end
			end
			3269: begin
				if(in == 0) begin
					state<=3270;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=7159;
					out<=219;
				end
				if(in == 3) begin
					state<=1338;
					out<=220;
				end
				if(in == 4) begin
					state<=5227;
					out<=221;
				end
			end
			3270: begin
				if(in == 0) begin
					state<=3271;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=7160;
					out<=224;
				end
				if(in == 3) begin
					state<=1339;
					out<=225;
				end
				if(in == 4) begin
					state<=5228;
					out<=226;
				end
			end
			3271: begin
				if(in == 0) begin
					state<=3272;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=7161;
					out<=229;
				end
				if(in == 3) begin
					state<=1340;
					out<=230;
				end
				if(in == 4) begin
					state<=5229;
					out<=231;
				end
			end
			3272: begin
				if(in == 0) begin
					state<=3273;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=7162;
					out<=234;
				end
				if(in == 3) begin
					state<=1341;
					out<=235;
				end
				if(in == 4) begin
					state<=5230;
					out<=236;
				end
			end
			3273: begin
				if(in == 0) begin
					state<=3274;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=7163;
					out<=239;
				end
				if(in == 3) begin
					state<=1342;
					out<=240;
				end
				if(in == 4) begin
					state<=5231;
					out<=241;
				end
			end
			3274: begin
				if(in == 0) begin
					state<=3275;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=7164;
					out<=244;
				end
				if(in == 3) begin
					state<=1343;
					out<=245;
				end
				if(in == 4) begin
					state<=5232;
					out<=246;
				end
			end
			3275: begin
				if(in == 0) begin
					state<=3276;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=7165;
					out<=249;
				end
				if(in == 3) begin
					state<=1344;
					out<=250;
				end
				if(in == 4) begin
					state<=5233;
					out<=251;
				end
			end
			3276: begin
				if(in == 0) begin
					state<=3277;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=7166;
					out<=254;
				end
				if(in == 3) begin
					state<=1345;
					out<=255;
				end
				if(in == 4) begin
					state<=5234;
					out<=0;
				end
			end
			3277: begin
				if(in == 0) begin
					state<=3278;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=7167;
					out<=3;
				end
				if(in == 3) begin
					state<=1346;
					out<=4;
				end
				if(in == 4) begin
					state<=5235;
					out<=5;
				end
			end
			3278: begin
				if(in == 0) begin
					state<=3279;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=7168;
					out<=8;
				end
				if(in == 3) begin
					state<=1347;
					out<=9;
				end
				if(in == 4) begin
					state<=5236;
					out<=10;
				end
			end
			3279: begin
				if(in == 0) begin
					state<=3280;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=7169;
					out<=13;
				end
				if(in == 3) begin
					state<=1348;
					out<=14;
				end
				if(in == 4) begin
					state<=5237;
					out<=15;
				end
			end
			3280: begin
				if(in == 0) begin
					state<=3281;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=7170;
					out<=18;
				end
				if(in == 3) begin
					state<=1349;
					out<=19;
				end
				if(in == 4) begin
					state<=5238;
					out<=20;
				end
			end
			3281: begin
				if(in == 0) begin
					state<=3282;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=7171;
					out<=23;
				end
				if(in == 3) begin
					state<=1350;
					out<=24;
				end
				if(in == 4) begin
					state<=5239;
					out<=25;
				end
			end
			3282: begin
				if(in == 0) begin
					state<=3283;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=7172;
					out<=28;
				end
				if(in == 3) begin
					state<=1351;
					out<=29;
				end
				if(in == 4) begin
					state<=5240;
					out<=30;
				end
			end
			3283: begin
				if(in == 0) begin
					state<=3284;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=7173;
					out<=33;
				end
				if(in == 3) begin
					state<=1352;
					out<=34;
				end
				if(in == 4) begin
					state<=5241;
					out<=35;
				end
			end
			3284: begin
				if(in == 0) begin
					state<=3285;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=7174;
					out<=38;
				end
				if(in == 3) begin
					state<=1353;
					out<=39;
				end
				if(in == 4) begin
					state<=5242;
					out<=40;
				end
			end
			3285: begin
				if(in == 0) begin
					state<=3286;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=7175;
					out<=43;
				end
				if(in == 3) begin
					state<=1354;
					out<=44;
				end
				if(in == 4) begin
					state<=5243;
					out<=45;
				end
			end
			3286: begin
				if(in == 0) begin
					state<=3287;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=7176;
					out<=48;
				end
				if(in == 3) begin
					state<=1355;
					out<=49;
				end
				if(in == 4) begin
					state<=5244;
					out<=50;
				end
			end
			3287: begin
				if(in == 0) begin
					state<=3288;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=7177;
					out<=53;
				end
				if(in == 3) begin
					state<=1356;
					out<=54;
				end
				if(in == 4) begin
					state<=5245;
					out<=55;
				end
			end
			3288: begin
				if(in == 0) begin
					state<=3289;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=7178;
					out<=58;
				end
				if(in == 3) begin
					state<=1357;
					out<=59;
				end
				if(in == 4) begin
					state<=5246;
					out<=60;
				end
			end
			3289: begin
				if(in == 0) begin
					state<=3290;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=7179;
					out<=63;
				end
				if(in == 3) begin
					state<=1358;
					out<=64;
				end
				if(in == 4) begin
					state<=5247;
					out<=65;
				end
			end
			3290: begin
				if(in == 0) begin
					state<=3291;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=7180;
					out<=68;
				end
				if(in == 3) begin
					state<=1359;
					out<=69;
				end
				if(in == 4) begin
					state<=5248;
					out<=70;
				end
			end
			3291: begin
				if(in == 0) begin
					state<=2049;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=5938;
					out<=73;
				end
				if(in == 3) begin
					state<=51;
					out<=74;
				end
				if(in == 4) begin
					state<=3949;
					out<=75;
				end
			end
			3292: begin
				if(in == 0) begin
					state<=3293;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=7182;
					out<=78;
				end
				if(in == 3) begin
					state<=1361;
					out<=79;
				end
				if(in == 4) begin
					state<=5250;
					out<=80;
				end
			end
			3293: begin
				if(in == 0) begin
					state<=3294;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=7183;
					out<=83;
				end
				if(in == 3) begin
					state<=1362;
					out<=84;
				end
				if(in == 4) begin
					state<=5251;
					out<=85;
				end
			end
			3294: begin
				if(in == 0) begin
					state<=3295;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=7184;
					out<=88;
				end
				if(in == 3) begin
					state<=1363;
					out<=89;
				end
				if(in == 4) begin
					state<=5252;
					out<=90;
				end
			end
			3295: begin
				if(in == 0) begin
					state<=3296;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=7185;
					out<=93;
				end
				if(in == 3) begin
					state<=1364;
					out<=94;
				end
				if(in == 4) begin
					state<=5253;
					out<=95;
				end
			end
			3296: begin
				if(in == 0) begin
					state<=3297;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=7186;
					out<=98;
				end
				if(in == 3) begin
					state<=1365;
					out<=99;
				end
				if(in == 4) begin
					state<=5254;
					out<=100;
				end
			end
			3297: begin
				if(in == 0) begin
					state<=3298;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=7187;
					out<=103;
				end
				if(in == 3) begin
					state<=1366;
					out<=104;
				end
				if(in == 4) begin
					state<=5255;
					out<=105;
				end
			end
			3298: begin
				if(in == 0) begin
					state<=3299;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=7188;
					out<=108;
				end
				if(in == 3) begin
					state<=1367;
					out<=109;
				end
				if(in == 4) begin
					state<=5256;
					out<=110;
				end
			end
			3299: begin
				if(in == 0) begin
					state<=3300;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=7189;
					out<=113;
				end
				if(in == 3) begin
					state<=1368;
					out<=114;
				end
				if(in == 4) begin
					state<=5257;
					out<=115;
				end
			end
			3300: begin
				if(in == 0) begin
					state<=3301;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=7190;
					out<=118;
				end
				if(in == 3) begin
					state<=1369;
					out<=119;
				end
				if(in == 4) begin
					state<=5258;
					out<=120;
				end
			end
			3301: begin
				if(in == 0) begin
					state<=3302;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=7191;
					out<=123;
				end
				if(in == 3) begin
					state<=1370;
					out<=124;
				end
				if(in == 4) begin
					state<=5259;
					out<=125;
				end
			end
			3302: begin
				if(in == 0) begin
					state<=3303;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=7192;
					out<=128;
				end
				if(in == 3) begin
					state<=1371;
					out<=129;
				end
				if(in == 4) begin
					state<=5260;
					out<=130;
				end
			end
			3303: begin
				if(in == 0) begin
					state<=3304;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=7193;
					out<=133;
				end
				if(in == 3) begin
					state<=1372;
					out<=134;
				end
				if(in == 4) begin
					state<=5261;
					out<=135;
				end
			end
			3304: begin
				if(in == 0) begin
					state<=3305;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=7194;
					out<=138;
				end
				if(in == 3) begin
					state<=1373;
					out<=139;
				end
				if(in == 4) begin
					state<=5262;
					out<=140;
				end
			end
			3305: begin
				if(in == 0) begin
					state<=3306;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=7195;
					out<=143;
				end
				if(in == 3) begin
					state<=1374;
					out<=144;
				end
				if(in == 4) begin
					state<=5263;
					out<=145;
				end
			end
			3306: begin
				if(in == 0) begin
					state<=3307;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=7196;
					out<=148;
				end
				if(in == 3) begin
					state<=1375;
					out<=149;
				end
				if(in == 4) begin
					state<=5264;
					out<=150;
				end
			end
			3307: begin
				if(in == 0) begin
					state<=3308;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=7197;
					out<=153;
				end
				if(in == 3) begin
					state<=1376;
					out<=154;
				end
				if(in == 4) begin
					state<=5265;
					out<=155;
				end
			end
			3308: begin
				if(in == 0) begin
					state<=3309;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=7198;
					out<=158;
				end
				if(in == 3) begin
					state<=1377;
					out<=159;
				end
				if(in == 4) begin
					state<=5266;
					out<=160;
				end
			end
			3309: begin
				if(in == 0) begin
					state<=3310;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=7199;
					out<=163;
				end
				if(in == 3) begin
					state<=1378;
					out<=164;
				end
				if(in == 4) begin
					state<=5267;
					out<=165;
				end
			end
			3310: begin
				if(in == 0) begin
					state<=3311;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=7200;
					out<=168;
				end
				if(in == 3) begin
					state<=1379;
					out<=169;
				end
				if(in == 4) begin
					state<=5268;
					out<=170;
				end
			end
			3311: begin
				if(in == 0) begin
					state<=3312;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=7201;
					out<=173;
				end
				if(in == 3) begin
					state<=1380;
					out<=174;
				end
				if(in == 4) begin
					state<=5269;
					out<=175;
				end
			end
			3312: begin
				if(in == 0) begin
					state<=3313;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=7202;
					out<=178;
				end
				if(in == 3) begin
					state<=1381;
					out<=179;
				end
				if(in == 4) begin
					state<=5270;
					out<=180;
				end
			end
			3313: begin
				if(in == 0) begin
					state<=3314;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=7203;
					out<=183;
				end
				if(in == 3) begin
					state<=1382;
					out<=184;
				end
				if(in == 4) begin
					state<=5271;
					out<=185;
				end
			end
			3314: begin
				if(in == 0) begin
					state<=3315;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=7204;
					out<=188;
				end
				if(in == 3) begin
					state<=1383;
					out<=189;
				end
				if(in == 4) begin
					state<=5272;
					out<=190;
				end
			end
			3315: begin
				if(in == 0) begin
					state<=3316;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=7205;
					out<=193;
				end
				if(in == 3) begin
					state<=1384;
					out<=194;
				end
				if(in == 4) begin
					state<=5273;
					out<=195;
				end
			end
			3316: begin
				if(in == 0) begin
					state<=3317;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=7206;
					out<=198;
				end
				if(in == 3) begin
					state<=1385;
					out<=199;
				end
				if(in == 4) begin
					state<=5274;
					out<=200;
				end
			end
			3317: begin
				if(in == 0) begin
					state<=3318;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=7207;
					out<=203;
				end
				if(in == 3) begin
					state<=1386;
					out<=204;
				end
				if(in == 4) begin
					state<=5275;
					out<=205;
				end
			end
			3318: begin
				if(in == 0) begin
					state<=3319;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=7208;
					out<=208;
				end
				if(in == 3) begin
					state<=1387;
					out<=209;
				end
				if(in == 4) begin
					state<=5276;
					out<=210;
				end
			end
			3319: begin
				if(in == 0) begin
					state<=3320;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=7209;
					out<=213;
				end
				if(in == 3) begin
					state<=1388;
					out<=214;
				end
				if(in == 4) begin
					state<=5277;
					out<=215;
				end
			end
			3320: begin
				if(in == 0) begin
					state<=3321;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=7210;
					out<=218;
				end
				if(in == 3) begin
					state<=1389;
					out<=219;
				end
				if(in == 4) begin
					state<=5278;
					out<=220;
				end
			end
			3321: begin
				if(in == 0) begin
					state<=3322;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=7211;
					out<=223;
				end
				if(in == 3) begin
					state<=1390;
					out<=224;
				end
				if(in == 4) begin
					state<=5279;
					out<=225;
				end
			end
			3322: begin
				if(in == 0) begin
					state<=2118;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=6007;
					out<=228;
				end
				if(in == 3) begin
					state<=120;
					out<=229;
				end
				if(in == 4) begin
					state<=4018;
					out<=230;
				end
			end
			3323: begin
				if(in == 0) begin
					state<=3324;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=7213;
					out<=233;
				end
				if(in == 3) begin
					state<=1392;
					out<=234;
				end
				if(in == 4) begin
					state<=5281;
					out<=235;
				end
			end
			3324: begin
				if(in == 0) begin
					state<=3325;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=7214;
					out<=238;
				end
				if(in == 3) begin
					state<=1393;
					out<=239;
				end
				if(in == 4) begin
					state<=5282;
					out<=240;
				end
			end
			3325: begin
				if(in == 0) begin
					state<=3326;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=7215;
					out<=243;
				end
				if(in == 3) begin
					state<=1394;
					out<=244;
				end
				if(in == 4) begin
					state<=5283;
					out<=245;
				end
			end
			3326: begin
				if(in == 0) begin
					state<=3327;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=7216;
					out<=248;
				end
				if(in == 3) begin
					state<=1395;
					out<=249;
				end
				if(in == 4) begin
					state<=5284;
					out<=250;
				end
			end
			3327: begin
				if(in == 0) begin
					state<=3328;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=7217;
					out<=253;
				end
				if(in == 3) begin
					state<=1396;
					out<=254;
				end
				if(in == 4) begin
					state<=5285;
					out<=255;
				end
			end
			3328: begin
				if(in == 0) begin
					state<=3329;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=7218;
					out<=2;
				end
				if(in == 3) begin
					state<=1397;
					out<=3;
				end
				if(in == 4) begin
					state<=5286;
					out<=4;
				end
			end
			3329: begin
				if(in == 0) begin
					state<=3330;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=7219;
					out<=7;
				end
				if(in == 3) begin
					state<=1398;
					out<=8;
				end
				if(in == 4) begin
					state<=5287;
					out<=9;
				end
			end
			3330: begin
				if(in == 0) begin
					state<=3331;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=7220;
					out<=12;
				end
				if(in == 3) begin
					state<=1399;
					out<=13;
				end
				if(in == 4) begin
					state<=5288;
					out<=14;
				end
			end
			3331: begin
				if(in == 0) begin
					state<=3332;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=7221;
					out<=17;
				end
				if(in == 3) begin
					state<=1400;
					out<=18;
				end
				if(in == 4) begin
					state<=5289;
					out<=19;
				end
			end
			3332: begin
				if(in == 0) begin
					state<=3333;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=7222;
					out<=22;
				end
				if(in == 3) begin
					state<=1401;
					out<=23;
				end
				if(in == 4) begin
					state<=5290;
					out<=24;
				end
			end
			3333: begin
				if(in == 0) begin
					state<=3334;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=7223;
					out<=27;
				end
				if(in == 3) begin
					state<=1402;
					out<=28;
				end
				if(in == 4) begin
					state<=5291;
					out<=29;
				end
			end
			3334: begin
				if(in == 0) begin
					state<=3335;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=7224;
					out<=32;
				end
				if(in == 3) begin
					state<=1403;
					out<=33;
				end
				if(in == 4) begin
					state<=5292;
					out<=34;
				end
			end
			3335: begin
				if(in == 0) begin
					state<=3336;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=7225;
					out<=37;
				end
				if(in == 3) begin
					state<=1404;
					out<=38;
				end
				if(in == 4) begin
					state<=5293;
					out<=39;
				end
			end
			3336: begin
				if(in == 0) begin
					state<=3337;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=7226;
					out<=42;
				end
				if(in == 3) begin
					state<=1405;
					out<=43;
				end
				if(in == 4) begin
					state<=5294;
					out<=44;
				end
			end
			3337: begin
				if(in == 0) begin
					state<=3338;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=7227;
					out<=47;
				end
				if(in == 3) begin
					state<=1406;
					out<=48;
				end
				if(in == 4) begin
					state<=5295;
					out<=49;
				end
			end
			3338: begin
				if(in == 0) begin
					state<=3339;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=7228;
					out<=52;
				end
				if(in == 3) begin
					state<=1407;
					out<=53;
				end
				if(in == 4) begin
					state<=5296;
					out<=54;
				end
			end
			3339: begin
				if(in == 0) begin
					state<=3340;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=7229;
					out<=57;
				end
				if(in == 3) begin
					state<=1408;
					out<=58;
				end
				if(in == 4) begin
					state<=5297;
					out<=59;
				end
			end
			3340: begin
				if(in == 0) begin
					state<=3341;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=7230;
					out<=62;
				end
				if(in == 3) begin
					state<=1409;
					out<=63;
				end
				if(in == 4) begin
					state<=5298;
					out<=64;
				end
			end
			3341: begin
				if(in == 0) begin
					state<=3342;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=7231;
					out<=67;
				end
				if(in == 3) begin
					state<=1410;
					out<=68;
				end
				if(in == 4) begin
					state<=5299;
					out<=69;
				end
			end
			3342: begin
				if(in == 0) begin
					state<=3343;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=7232;
					out<=72;
				end
				if(in == 3) begin
					state<=1411;
					out<=73;
				end
				if(in == 4) begin
					state<=5300;
					out<=74;
				end
			end
			3343: begin
				if(in == 0) begin
					state<=3344;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=7233;
					out<=77;
				end
				if(in == 3) begin
					state<=1412;
					out<=78;
				end
				if(in == 4) begin
					state<=5301;
					out<=79;
				end
			end
			3344: begin
				if(in == 0) begin
					state<=3345;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=7234;
					out<=82;
				end
				if(in == 3) begin
					state<=1413;
					out<=83;
				end
				if(in == 4) begin
					state<=5302;
					out<=84;
				end
			end
			3345: begin
				if(in == 0) begin
					state<=3346;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=7235;
					out<=87;
				end
				if(in == 3) begin
					state<=1414;
					out<=88;
				end
				if(in == 4) begin
					state<=5303;
					out<=89;
				end
			end
			3346: begin
				if(in == 0) begin
					state<=3347;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=7236;
					out<=92;
				end
				if(in == 3) begin
					state<=1415;
					out<=93;
				end
				if(in == 4) begin
					state<=5304;
					out<=94;
				end
			end
			3347: begin
				if(in == 0) begin
					state<=3348;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=7237;
					out<=97;
				end
				if(in == 3) begin
					state<=1416;
					out<=98;
				end
				if(in == 4) begin
					state<=5305;
					out<=99;
				end
			end
			3348: begin
				if(in == 0) begin
					state<=3349;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=7238;
					out<=102;
				end
				if(in == 3) begin
					state<=1417;
					out<=103;
				end
				if(in == 4) begin
					state<=5306;
					out<=104;
				end
			end
			3349: begin
				if(in == 0) begin
					state<=3350;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=7239;
					out<=107;
				end
				if(in == 3) begin
					state<=1418;
					out<=108;
				end
				if(in == 4) begin
					state<=5307;
					out<=109;
				end
			end
			3350: begin
				if(in == 0) begin
					state<=3351;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=7240;
					out<=112;
				end
				if(in == 3) begin
					state<=1419;
					out<=113;
				end
				if(in == 4) begin
					state<=5308;
					out<=114;
				end
			end
			3351: begin
				if(in == 0) begin
					state<=3352;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=7241;
					out<=117;
				end
				if(in == 3) begin
					state<=1420;
					out<=118;
				end
				if(in == 4) begin
					state<=5309;
					out<=119;
				end
			end
			3352: begin
				if(in == 0) begin
					state<=3353;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=7242;
					out<=122;
				end
				if(in == 3) begin
					state<=1421;
					out<=123;
				end
				if(in == 4) begin
					state<=5310;
					out<=124;
				end
			end
			3353: begin
				if(in == 0) begin
					state<=2187;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=6076;
					out<=127;
				end
				if(in == 3) begin
					state<=189;
					out<=128;
				end
				if(in == 4) begin
					state<=4087;
					out<=129;
				end
			end
			3354: begin
				if(in == 0) begin
					state<=3355;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=7244;
					out<=132;
				end
				if(in == 3) begin
					state<=1423;
					out<=133;
				end
				if(in == 4) begin
					state<=5312;
					out<=134;
				end
			end
			3355: begin
				if(in == 0) begin
					state<=3356;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=7245;
					out<=137;
				end
				if(in == 3) begin
					state<=1424;
					out<=138;
				end
				if(in == 4) begin
					state<=5313;
					out<=139;
				end
			end
			3356: begin
				if(in == 0) begin
					state<=3357;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=7246;
					out<=142;
				end
				if(in == 3) begin
					state<=1425;
					out<=143;
				end
				if(in == 4) begin
					state<=5314;
					out<=144;
				end
			end
			3357: begin
				if(in == 0) begin
					state<=3358;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=7247;
					out<=147;
				end
				if(in == 3) begin
					state<=1426;
					out<=148;
				end
				if(in == 4) begin
					state<=5315;
					out<=149;
				end
			end
			3358: begin
				if(in == 0) begin
					state<=3359;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=7248;
					out<=152;
				end
				if(in == 3) begin
					state<=1427;
					out<=153;
				end
				if(in == 4) begin
					state<=5316;
					out<=154;
				end
			end
			3359: begin
				if(in == 0) begin
					state<=3360;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=7249;
					out<=157;
				end
				if(in == 3) begin
					state<=1428;
					out<=158;
				end
				if(in == 4) begin
					state<=5317;
					out<=159;
				end
			end
			3360: begin
				if(in == 0) begin
					state<=3361;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=7250;
					out<=162;
				end
				if(in == 3) begin
					state<=1429;
					out<=163;
				end
				if(in == 4) begin
					state<=5318;
					out<=164;
				end
			end
			3361: begin
				if(in == 0) begin
					state<=3362;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=7251;
					out<=167;
				end
				if(in == 3) begin
					state<=1430;
					out<=168;
				end
				if(in == 4) begin
					state<=5319;
					out<=169;
				end
			end
			3362: begin
				if(in == 0) begin
					state<=3363;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=7252;
					out<=172;
				end
				if(in == 3) begin
					state<=1431;
					out<=173;
				end
				if(in == 4) begin
					state<=5320;
					out<=174;
				end
			end
			3363: begin
				if(in == 0) begin
					state<=3364;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=7253;
					out<=177;
				end
				if(in == 3) begin
					state<=1432;
					out<=178;
				end
				if(in == 4) begin
					state<=5321;
					out<=179;
				end
			end
			3364: begin
				if(in == 0) begin
					state<=3365;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=7254;
					out<=182;
				end
				if(in == 3) begin
					state<=1433;
					out<=183;
				end
				if(in == 4) begin
					state<=5322;
					out<=184;
				end
			end
			3365: begin
				if(in == 0) begin
					state<=3366;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=7255;
					out<=187;
				end
				if(in == 3) begin
					state<=1434;
					out<=188;
				end
				if(in == 4) begin
					state<=5323;
					out<=189;
				end
			end
			3366: begin
				if(in == 0) begin
					state<=3367;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=7256;
					out<=192;
				end
				if(in == 3) begin
					state<=1435;
					out<=193;
				end
				if(in == 4) begin
					state<=5324;
					out<=194;
				end
			end
			3367: begin
				if(in == 0) begin
					state<=3368;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=7257;
					out<=197;
				end
				if(in == 3) begin
					state<=1436;
					out<=198;
				end
				if(in == 4) begin
					state<=5325;
					out<=199;
				end
			end
			3368: begin
				if(in == 0) begin
					state<=3369;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=7258;
					out<=202;
				end
				if(in == 3) begin
					state<=1437;
					out<=203;
				end
				if(in == 4) begin
					state<=5326;
					out<=204;
				end
			end
			3369: begin
				if(in == 0) begin
					state<=3370;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=7259;
					out<=207;
				end
				if(in == 3) begin
					state<=1438;
					out<=208;
				end
				if(in == 4) begin
					state<=5327;
					out<=209;
				end
			end
			3370: begin
				if(in == 0) begin
					state<=3371;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=7260;
					out<=212;
				end
				if(in == 3) begin
					state<=1439;
					out<=213;
				end
				if(in == 4) begin
					state<=5328;
					out<=214;
				end
			end
			3371: begin
				if(in == 0) begin
					state<=3372;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=7261;
					out<=217;
				end
				if(in == 3) begin
					state<=1440;
					out<=218;
				end
				if(in == 4) begin
					state<=5329;
					out<=219;
				end
			end
			3372: begin
				if(in == 0) begin
					state<=3373;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=7262;
					out<=222;
				end
				if(in == 3) begin
					state<=1441;
					out<=223;
				end
				if(in == 4) begin
					state<=5330;
					out<=224;
				end
			end
			3373: begin
				if(in == 0) begin
					state<=3374;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=7263;
					out<=227;
				end
				if(in == 3) begin
					state<=1442;
					out<=228;
				end
				if(in == 4) begin
					state<=5331;
					out<=229;
				end
			end
			3374: begin
				if(in == 0) begin
					state<=3375;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=7264;
					out<=232;
				end
				if(in == 3) begin
					state<=1443;
					out<=233;
				end
				if(in == 4) begin
					state<=5332;
					out<=234;
				end
			end
			3375: begin
				if(in == 0) begin
					state<=3376;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=7265;
					out<=237;
				end
				if(in == 3) begin
					state<=1444;
					out<=238;
				end
				if(in == 4) begin
					state<=5333;
					out<=239;
				end
			end
			3376: begin
				if(in == 0) begin
					state<=3377;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=7266;
					out<=242;
				end
				if(in == 3) begin
					state<=1445;
					out<=243;
				end
				if(in == 4) begin
					state<=5334;
					out<=244;
				end
			end
			3377: begin
				if(in == 0) begin
					state<=3378;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=7267;
					out<=247;
				end
				if(in == 3) begin
					state<=1446;
					out<=248;
				end
				if(in == 4) begin
					state<=5335;
					out<=249;
				end
			end
			3378: begin
				if(in == 0) begin
					state<=3379;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=7268;
					out<=252;
				end
				if(in == 3) begin
					state<=1447;
					out<=253;
				end
				if(in == 4) begin
					state<=5336;
					out<=254;
				end
			end
			3379: begin
				if(in == 0) begin
					state<=3380;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=7269;
					out<=1;
				end
				if(in == 3) begin
					state<=1448;
					out<=2;
				end
				if(in == 4) begin
					state<=5337;
					out<=3;
				end
			end
			3380: begin
				if(in == 0) begin
					state<=3381;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=7270;
					out<=6;
				end
				if(in == 3) begin
					state<=1449;
					out<=7;
				end
				if(in == 4) begin
					state<=5338;
					out<=8;
				end
			end
			3381: begin
				if(in == 0) begin
					state<=3382;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=7271;
					out<=11;
				end
				if(in == 3) begin
					state<=1450;
					out<=12;
				end
				if(in == 4) begin
					state<=5339;
					out<=13;
				end
			end
			3382: begin
				if(in == 0) begin
					state<=3383;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=7272;
					out<=16;
				end
				if(in == 3) begin
					state<=1451;
					out<=17;
				end
				if(in == 4) begin
					state<=5340;
					out<=18;
				end
			end
			3383: begin
				if(in == 0) begin
					state<=3384;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=7273;
					out<=21;
				end
				if(in == 3) begin
					state<=1452;
					out<=22;
				end
				if(in == 4) begin
					state<=5341;
					out<=23;
				end
			end
			3384: begin
				if(in == 0) begin
					state<=2256;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=6145;
					out<=26;
				end
				if(in == 3) begin
					state<=258;
					out<=27;
				end
				if(in == 4) begin
					state<=4156;
					out<=28;
				end
			end
			3385: begin
				if(in == 0) begin
					state<=3386;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=7275;
					out<=31;
				end
				if(in == 3) begin
					state<=1000;
					out<=32;
				end
				if(in == 4) begin
					state<=4898;
					out<=33;
				end
			end
			3386: begin
				if(in == 0) begin
					state<=3387;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=7276;
					out<=36;
				end
				if(in == 3) begin
					state<=1001;
					out<=37;
				end
				if(in == 4) begin
					state<=4899;
					out<=38;
				end
			end
			3387: begin
				if(in == 0) begin
					state<=3388;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=7277;
					out<=41;
				end
				if(in == 3) begin
					state<=1002;
					out<=42;
				end
				if(in == 4) begin
					state<=4900;
					out<=43;
				end
			end
			3388: begin
				if(in == 0) begin
					state<=3389;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=7278;
					out<=46;
				end
				if(in == 3) begin
					state<=1003;
					out<=47;
				end
				if(in == 4) begin
					state<=4901;
					out<=48;
				end
			end
			3389: begin
				if(in == 0) begin
					state<=3390;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=7279;
					out<=51;
				end
				if(in == 3) begin
					state<=1004;
					out<=52;
				end
				if(in == 4) begin
					state<=4902;
					out<=53;
				end
			end
			3390: begin
				if(in == 0) begin
					state<=3391;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=7280;
					out<=56;
				end
				if(in == 3) begin
					state<=1005;
					out<=57;
				end
				if(in == 4) begin
					state<=4903;
					out<=58;
				end
			end
			3391: begin
				if(in == 0) begin
					state<=3392;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=7281;
					out<=61;
				end
				if(in == 3) begin
					state<=1006;
					out<=62;
				end
				if(in == 4) begin
					state<=4904;
					out<=63;
				end
			end
			3392: begin
				if(in == 0) begin
					state<=3393;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=7282;
					out<=66;
				end
				if(in == 3) begin
					state<=1007;
					out<=67;
				end
				if(in == 4) begin
					state<=4905;
					out<=68;
				end
			end
			3393: begin
				if(in == 0) begin
					state<=3394;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=7283;
					out<=71;
				end
				if(in == 3) begin
					state<=1008;
					out<=72;
				end
				if(in == 4) begin
					state<=4906;
					out<=73;
				end
			end
			3394: begin
				if(in == 0) begin
					state<=3395;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=7284;
					out<=76;
				end
				if(in == 3) begin
					state<=1009;
					out<=77;
				end
				if(in == 4) begin
					state<=4907;
					out<=78;
				end
			end
			3395: begin
				if(in == 0) begin
					state<=3396;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=7285;
					out<=81;
				end
				if(in == 3) begin
					state<=1010;
					out<=82;
				end
				if(in == 4) begin
					state<=4908;
					out<=83;
				end
			end
			3396: begin
				if(in == 0) begin
					state<=3397;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=7286;
					out<=86;
				end
				if(in == 3) begin
					state<=1011;
					out<=87;
				end
				if(in == 4) begin
					state<=4909;
					out<=88;
				end
			end
			3397: begin
				if(in == 0) begin
					state<=3398;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=7287;
					out<=91;
				end
				if(in == 3) begin
					state<=1012;
					out<=92;
				end
				if(in == 4) begin
					state<=4910;
					out<=93;
				end
			end
			3398: begin
				if(in == 0) begin
					state<=3399;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=7288;
					out<=96;
				end
				if(in == 3) begin
					state<=1013;
					out<=97;
				end
				if(in == 4) begin
					state<=4911;
					out<=98;
				end
			end
			3399: begin
				if(in == 0) begin
					state<=3400;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=7289;
					out<=101;
				end
				if(in == 3) begin
					state<=1014;
					out<=102;
				end
				if(in == 4) begin
					state<=4912;
					out<=103;
				end
			end
			3400: begin
				if(in == 0) begin
					state<=3401;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=7290;
					out<=106;
				end
				if(in == 3) begin
					state<=1015;
					out<=107;
				end
				if(in == 4) begin
					state<=4913;
					out<=108;
				end
			end
			3401: begin
				if(in == 0) begin
					state<=3402;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=7291;
					out<=111;
				end
				if(in == 3) begin
					state<=1016;
					out<=112;
				end
				if(in == 4) begin
					state<=4914;
					out<=113;
				end
			end
			3402: begin
				if(in == 0) begin
					state<=3403;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=7292;
					out<=116;
				end
				if(in == 3) begin
					state<=1017;
					out<=117;
				end
				if(in == 4) begin
					state<=4915;
					out<=118;
				end
			end
			3403: begin
				if(in == 0) begin
					state<=3404;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=7293;
					out<=121;
				end
				if(in == 3) begin
					state<=1018;
					out<=122;
				end
				if(in == 4) begin
					state<=4916;
					out<=123;
				end
			end
			3404: begin
				if(in == 0) begin
					state<=3405;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=7294;
					out<=126;
				end
				if(in == 3) begin
					state<=1019;
					out<=127;
				end
				if(in == 4) begin
					state<=4917;
					out<=128;
				end
			end
			3405: begin
				if(in == 0) begin
					state<=3406;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=7295;
					out<=131;
				end
				if(in == 3) begin
					state<=1020;
					out<=132;
				end
				if(in == 4) begin
					state<=4918;
					out<=133;
				end
			end
			3406: begin
				if(in == 0) begin
					state<=3407;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=7296;
					out<=136;
				end
				if(in == 3) begin
					state<=1021;
					out<=137;
				end
				if(in == 4) begin
					state<=4919;
					out<=138;
				end
			end
			3407: begin
				if(in == 0) begin
					state<=3408;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=7297;
					out<=141;
				end
				if(in == 3) begin
					state<=1022;
					out<=142;
				end
				if(in == 4) begin
					state<=4920;
					out<=143;
				end
			end
			3408: begin
				if(in == 0) begin
					state<=3409;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=7298;
					out<=146;
				end
				if(in == 3) begin
					state<=1023;
					out<=147;
				end
				if(in == 4) begin
					state<=4921;
					out<=148;
				end
			end
			3409: begin
				if(in == 0) begin
					state<=3410;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=7299;
					out<=151;
				end
				if(in == 3) begin
					state<=1024;
					out<=152;
				end
				if(in == 4) begin
					state<=4922;
					out<=153;
				end
			end
			3410: begin
				if(in == 0) begin
					state<=3411;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=7300;
					out<=156;
				end
				if(in == 3) begin
					state<=1025;
					out<=157;
				end
				if(in == 4) begin
					state<=4923;
					out<=158;
				end
			end
			3411: begin
				if(in == 0) begin
					state<=3412;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=7301;
					out<=161;
				end
				if(in == 3) begin
					state<=1026;
					out<=162;
				end
				if(in == 4) begin
					state<=4924;
					out<=163;
				end
			end
			3412: begin
				if(in == 0) begin
					state<=3413;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=7302;
					out<=166;
				end
				if(in == 3) begin
					state<=1027;
					out<=167;
				end
				if(in == 4) begin
					state<=4925;
					out<=168;
				end
			end
			3413: begin
				if(in == 0) begin
					state<=3414;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=7303;
					out<=171;
				end
				if(in == 3) begin
					state<=1028;
					out<=172;
				end
				if(in == 4) begin
					state<=4926;
					out<=173;
				end
			end
			3414: begin
				if(in == 0) begin
					state<=3415;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=7304;
					out<=176;
				end
				if(in == 3) begin
					state<=1029;
					out<=177;
				end
				if(in == 4) begin
					state<=4927;
					out<=178;
				end
			end
			3415: begin
				if(in == 0) begin
					state<=2394;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=6283;
					out<=181;
				end
				if(in == 3) begin
					state<=396;
					out<=182;
				end
				if(in == 4) begin
					state<=4294;
					out<=183;
				end
			end
			3416: begin
				if(in == 0) begin
					state<=3417;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=7306;
					out<=186;
				end
				if(in == 3) begin
					state<=1485;
					out<=187;
				end
				if(in == 4) begin
					state<=5374;
					out<=188;
				end
			end
			3417: begin
				if(in == 0) begin
					state<=3418;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=7307;
					out<=191;
				end
				if(in == 3) begin
					state<=1486;
					out<=192;
				end
				if(in == 4) begin
					state<=5375;
					out<=193;
				end
			end
			3418: begin
				if(in == 0) begin
					state<=3419;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=7308;
					out<=196;
				end
				if(in == 3) begin
					state<=1487;
					out<=197;
				end
				if(in == 4) begin
					state<=5376;
					out<=198;
				end
			end
			3419: begin
				if(in == 0) begin
					state<=3420;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=7309;
					out<=201;
				end
				if(in == 3) begin
					state<=1488;
					out<=202;
				end
				if(in == 4) begin
					state<=5377;
					out<=203;
				end
			end
			3420: begin
				if(in == 0) begin
					state<=3421;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=7310;
					out<=206;
				end
				if(in == 3) begin
					state<=1489;
					out<=207;
				end
				if(in == 4) begin
					state<=5378;
					out<=208;
				end
			end
			3421: begin
				if(in == 0) begin
					state<=3422;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=7311;
					out<=211;
				end
				if(in == 3) begin
					state<=1490;
					out<=212;
				end
				if(in == 4) begin
					state<=5379;
					out<=213;
				end
			end
			3422: begin
				if(in == 0) begin
					state<=3423;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=7312;
					out<=216;
				end
				if(in == 3) begin
					state<=1491;
					out<=217;
				end
				if(in == 4) begin
					state<=5380;
					out<=218;
				end
			end
			3423: begin
				if(in == 0) begin
					state<=3424;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=7313;
					out<=221;
				end
				if(in == 3) begin
					state<=1492;
					out<=222;
				end
				if(in == 4) begin
					state<=5381;
					out<=223;
				end
			end
			3424: begin
				if(in == 0) begin
					state<=3425;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=7314;
					out<=226;
				end
				if(in == 3) begin
					state<=1493;
					out<=227;
				end
				if(in == 4) begin
					state<=5382;
					out<=228;
				end
			end
			3425: begin
				if(in == 0) begin
					state<=3426;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=7315;
					out<=231;
				end
				if(in == 3) begin
					state<=1494;
					out<=232;
				end
				if(in == 4) begin
					state<=5383;
					out<=233;
				end
			end
			3426: begin
				if(in == 0) begin
					state<=3427;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=7316;
					out<=236;
				end
				if(in == 3) begin
					state<=1495;
					out<=237;
				end
				if(in == 4) begin
					state<=5384;
					out<=238;
				end
			end
			3427: begin
				if(in == 0) begin
					state<=3428;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=7317;
					out<=241;
				end
				if(in == 3) begin
					state<=1496;
					out<=242;
				end
				if(in == 4) begin
					state<=5385;
					out<=243;
				end
			end
			3428: begin
				if(in == 0) begin
					state<=3429;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=7318;
					out<=246;
				end
				if(in == 3) begin
					state<=1497;
					out<=247;
				end
				if(in == 4) begin
					state<=5386;
					out<=248;
				end
			end
			3429: begin
				if(in == 0) begin
					state<=3430;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=7319;
					out<=251;
				end
				if(in == 3) begin
					state<=1498;
					out<=252;
				end
				if(in == 4) begin
					state<=5387;
					out<=253;
				end
			end
			3430: begin
				if(in == 0) begin
					state<=3431;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=7320;
					out<=0;
				end
				if(in == 3) begin
					state<=1499;
					out<=1;
				end
				if(in == 4) begin
					state<=5388;
					out<=2;
				end
			end
			3431: begin
				if(in == 0) begin
					state<=3432;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=7321;
					out<=5;
				end
				if(in == 3) begin
					state<=1500;
					out<=6;
				end
				if(in == 4) begin
					state<=5389;
					out<=7;
				end
			end
			3432: begin
				if(in == 0) begin
					state<=3433;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=7322;
					out<=10;
				end
				if(in == 3) begin
					state<=1501;
					out<=11;
				end
				if(in == 4) begin
					state<=5390;
					out<=12;
				end
			end
			3433: begin
				if(in == 0) begin
					state<=3434;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=7323;
					out<=15;
				end
				if(in == 3) begin
					state<=1502;
					out<=16;
				end
				if(in == 4) begin
					state<=5391;
					out<=17;
				end
			end
			3434: begin
				if(in == 0) begin
					state<=3435;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=7324;
					out<=20;
				end
				if(in == 3) begin
					state<=1503;
					out<=21;
				end
				if(in == 4) begin
					state<=5392;
					out<=22;
				end
			end
			3435: begin
				if(in == 0) begin
					state<=3436;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=7325;
					out<=25;
				end
				if(in == 3) begin
					state<=1504;
					out<=26;
				end
				if(in == 4) begin
					state<=5393;
					out<=27;
				end
			end
			3436: begin
				if(in == 0) begin
					state<=3437;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=7326;
					out<=30;
				end
				if(in == 3) begin
					state<=1505;
					out<=31;
				end
				if(in == 4) begin
					state<=5394;
					out<=32;
				end
			end
			3437: begin
				if(in == 0) begin
					state<=3438;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=7327;
					out<=35;
				end
				if(in == 3) begin
					state<=1506;
					out<=36;
				end
				if(in == 4) begin
					state<=5395;
					out<=37;
				end
			end
			3438: begin
				if(in == 0) begin
					state<=3439;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=7328;
					out<=40;
				end
				if(in == 3) begin
					state<=1507;
					out<=41;
				end
				if(in == 4) begin
					state<=5396;
					out<=42;
				end
			end
			3439: begin
				if(in == 0) begin
					state<=3440;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=7329;
					out<=45;
				end
				if(in == 3) begin
					state<=1508;
					out<=46;
				end
				if(in == 4) begin
					state<=5397;
					out<=47;
				end
			end
			3440: begin
				if(in == 0) begin
					state<=3441;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=7330;
					out<=50;
				end
				if(in == 3) begin
					state<=1509;
					out<=51;
				end
				if(in == 4) begin
					state<=5398;
					out<=52;
				end
			end
			3441: begin
				if(in == 0) begin
					state<=3442;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=7331;
					out<=55;
				end
				if(in == 3) begin
					state<=1510;
					out<=56;
				end
				if(in == 4) begin
					state<=5399;
					out<=57;
				end
			end
			3442: begin
				if(in == 0) begin
					state<=3443;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=7332;
					out<=60;
				end
				if(in == 3) begin
					state<=1511;
					out<=61;
				end
				if(in == 4) begin
					state<=5400;
					out<=62;
				end
			end
			3443: begin
				if(in == 0) begin
					state<=3444;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=7333;
					out<=65;
				end
				if(in == 3) begin
					state<=1512;
					out<=66;
				end
				if(in == 4) begin
					state<=5401;
					out<=67;
				end
			end
			3444: begin
				if(in == 0) begin
					state<=3445;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=7334;
					out<=70;
				end
				if(in == 3) begin
					state<=1513;
					out<=71;
				end
				if(in == 4) begin
					state<=5402;
					out<=72;
				end
			end
			3445: begin
				if(in == 0) begin
					state<=3446;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=7335;
					out<=75;
				end
				if(in == 3) begin
					state<=1514;
					out<=76;
				end
				if(in == 4) begin
					state<=5403;
					out<=77;
				end
			end
			3446: begin
				if(in == 0) begin
					state<=2463;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=6352;
					out<=80;
				end
				if(in == 3) begin
					state<=465;
					out<=81;
				end
				if(in == 4) begin
					state<=4363;
					out<=82;
				end
			end
			3447: begin
				if(in == 0) begin
					state<=3448;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=7337;
					out<=85;
				end
				if(in == 3) begin
					state<=1516;
					out<=86;
				end
				if(in == 4) begin
					state<=5405;
					out<=87;
				end
			end
			3448: begin
				if(in == 0) begin
					state<=3449;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=7338;
					out<=90;
				end
				if(in == 3) begin
					state<=1517;
					out<=91;
				end
				if(in == 4) begin
					state<=5406;
					out<=92;
				end
			end
			3449: begin
				if(in == 0) begin
					state<=3450;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=7339;
					out<=95;
				end
				if(in == 3) begin
					state<=1518;
					out<=96;
				end
				if(in == 4) begin
					state<=5407;
					out<=97;
				end
			end
			3450: begin
				if(in == 0) begin
					state<=3451;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=7340;
					out<=100;
				end
				if(in == 3) begin
					state<=1519;
					out<=101;
				end
				if(in == 4) begin
					state<=5408;
					out<=102;
				end
			end
			3451: begin
				if(in == 0) begin
					state<=3452;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=7341;
					out<=105;
				end
				if(in == 3) begin
					state<=1520;
					out<=106;
				end
				if(in == 4) begin
					state<=5409;
					out<=107;
				end
			end
			3452: begin
				if(in == 0) begin
					state<=3453;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=7342;
					out<=110;
				end
				if(in == 3) begin
					state<=1521;
					out<=111;
				end
				if(in == 4) begin
					state<=5410;
					out<=112;
				end
			end
			3453: begin
				if(in == 0) begin
					state<=3454;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=7343;
					out<=115;
				end
				if(in == 3) begin
					state<=1522;
					out<=116;
				end
				if(in == 4) begin
					state<=5411;
					out<=117;
				end
			end
			3454: begin
				if(in == 0) begin
					state<=3455;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=7344;
					out<=120;
				end
				if(in == 3) begin
					state<=1523;
					out<=121;
				end
				if(in == 4) begin
					state<=5412;
					out<=122;
				end
			end
			3455: begin
				if(in == 0) begin
					state<=3456;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=7345;
					out<=125;
				end
				if(in == 3) begin
					state<=1524;
					out<=126;
				end
				if(in == 4) begin
					state<=5413;
					out<=127;
				end
			end
			3456: begin
				if(in == 0) begin
					state<=3457;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=7346;
					out<=130;
				end
				if(in == 3) begin
					state<=1525;
					out<=131;
				end
				if(in == 4) begin
					state<=5414;
					out<=132;
				end
			end
			3457: begin
				if(in == 0) begin
					state<=3458;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=7347;
					out<=135;
				end
				if(in == 3) begin
					state<=1526;
					out<=136;
				end
				if(in == 4) begin
					state<=5415;
					out<=137;
				end
			end
			3458: begin
				if(in == 0) begin
					state<=3459;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=7348;
					out<=140;
				end
				if(in == 3) begin
					state<=1527;
					out<=141;
				end
				if(in == 4) begin
					state<=5416;
					out<=142;
				end
			end
			3459: begin
				if(in == 0) begin
					state<=3460;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=7349;
					out<=145;
				end
				if(in == 3) begin
					state<=1528;
					out<=146;
				end
				if(in == 4) begin
					state<=5417;
					out<=147;
				end
			end
			3460: begin
				if(in == 0) begin
					state<=3461;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=7350;
					out<=150;
				end
				if(in == 3) begin
					state<=1529;
					out<=151;
				end
				if(in == 4) begin
					state<=5418;
					out<=152;
				end
			end
			3461: begin
				if(in == 0) begin
					state<=3462;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=7351;
					out<=155;
				end
				if(in == 3) begin
					state<=1530;
					out<=156;
				end
				if(in == 4) begin
					state<=5419;
					out<=157;
				end
			end
			3462: begin
				if(in == 0) begin
					state<=3463;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=7352;
					out<=160;
				end
				if(in == 3) begin
					state<=1531;
					out<=161;
				end
				if(in == 4) begin
					state<=5420;
					out<=162;
				end
			end
			3463: begin
				if(in == 0) begin
					state<=3464;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=7353;
					out<=165;
				end
				if(in == 3) begin
					state<=1532;
					out<=166;
				end
				if(in == 4) begin
					state<=5421;
					out<=167;
				end
			end
			3464: begin
				if(in == 0) begin
					state<=3465;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=7354;
					out<=170;
				end
				if(in == 3) begin
					state<=1533;
					out<=171;
				end
				if(in == 4) begin
					state<=5422;
					out<=172;
				end
			end
			3465: begin
				if(in == 0) begin
					state<=3466;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=7355;
					out<=175;
				end
				if(in == 3) begin
					state<=1534;
					out<=176;
				end
				if(in == 4) begin
					state<=5423;
					out<=177;
				end
			end
			3466: begin
				if(in == 0) begin
					state<=3467;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=7356;
					out<=180;
				end
				if(in == 3) begin
					state<=1535;
					out<=181;
				end
				if(in == 4) begin
					state<=5424;
					out<=182;
				end
			end
			3467: begin
				if(in == 0) begin
					state<=3468;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=7357;
					out<=185;
				end
				if(in == 3) begin
					state<=1536;
					out<=186;
				end
				if(in == 4) begin
					state<=5425;
					out<=187;
				end
			end
			3468: begin
				if(in == 0) begin
					state<=3469;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=7358;
					out<=190;
				end
				if(in == 3) begin
					state<=1537;
					out<=191;
				end
				if(in == 4) begin
					state<=5426;
					out<=192;
				end
			end
			3469: begin
				if(in == 0) begin
					state<=3470;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=7359;
					out<=195;
				end
				if(in == 3) begin
					state<=1538;
					out<=196;
				end
				if(in == 4) begin
					state<=5427;
					out<=197;
				end
			end
			3470: begin
				if(in == 0) begin
					state<=3471;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=7360;
					out<=200;
				end
				if(in == 3) begin
					state<=1539;
					out<=201;
				end
				if(in == 4) begin
					state<=5428;
					out<=202;
				end
			end
			3471: begin
				if(in == 0) begin
					state<=3472;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=7361;
					out<=205;
				end
				if(in == 3) begin
					state<=1540;
					out<=206;
				end
				if(in == 4) begin
					state<=5429;
					out<=207;
				end
			end
			3472: begin
				if(in == 0) begin
					state<=3473;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=7362;
					out<=210;
				end
				if(in == 3) begin
					state<=1541;
					out<=211;
				end
				if(in == 4) begin
					state<=5430;
					out<=212;
				end
			end
			3473: begin
				if(in == 0) begin
					state<=3474;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=7363;
					out<=215;
				end
				if(in == 3) begin
					state<=1542;
					out<=216;
				end
				if(in == 4) begin
					state<=5431;
					out<=217;
				end
			end
			3474: begin
				if(in == 0) begin
					state<=3475;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=7364;
					out<=220;
				end
				if(in == 3) begin
					state<=1543;
					out<=221;
				end
				if(in == 4) begin
					state<=5432;
					out<=222;
				end
			end
			3475: begin
				if(in == 0) begin
					state<=3476;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=7365;
					out<=225;
				end
				if(in == 3) begin
					state<=1544;
					out<=226;
				end
				if(in == 4) begin
					state<=5433;
					out<=227;
				end
			end
			3476: begin
				if(in == 0) begin
					state<=3477;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=7366;
					out<=230;
				end
				if(in == 3) begin
					state<=1545;
					out<=231;
				end
				if(in == 4) begin
					state<=5434;
					out<=232;
				end
			end
			3477: begin
				if(in == 0) begin
					state<=2532;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=6421;
					out<=235;
				end
				if(in == 3) begin
					state<=534;
					out<=236;
				end
				if(in == 4) begin
					state<=4432;
					out<=237;
				end
			end
			3478: begin
				if(in == 0) begin
					state<=3479;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=7368;
					out<=240;
				end
				if(in == 3) begin
					state<=1547;
					out<=241;
				end
				if(in == 4) begin
					state<=5436;
					out<=242;
				end
			end
			3479: begin
				if(in == 0) begin
					state<=3480;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=7369;
					out<=245;
				end
				if(in == 3) begin
					state<=1548;
					out<=246;
				end
				if(in == 4) begin
					state<=5437;
					out<=247;
				end
			end
			3480: begin
				if(in == 0) begin
					state<=3481;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=7370;
					out<=250;
				end
				if(in == 3) begin
					state<=1549;
					out<=251;
				end
				if(in == 4) begin
					state<=5438;
					out<=252;
				end
			end
			3481: begin
				if(in == 0) begin
					state<=3482;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=7371;
					out<=255;
				end
				if(in == 3) begin
					state<=1550;
					out<=0;
				end
				if(in == 4) begin
					state<=5439;
					out<=1;
				end
			end
			3482: begin
				if(in == 0) begin
					state<=3483;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=7372;
					out<=4;
				end
				if(in == 3) begin
					state<=1551;
					out<=5;
				end
				if(in == 4) begin
					state<=5440;
					out<=6;
				end
			end
			3483: begin
				if(in == 0) begin
					state<=3484;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=7373;
					out<=9;
				end
				if(in == 3) begin
					state<=1552;
					out<=10;
				end
				if(in == 4) begin
					state<=5441;
					out<=11;
				end
			end
			3484: begin
				if(in == 0) begin
					state<=3485;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=7374;
					out<=14;
				end
				if(in == 3) begin
					state<=1553;
					out<=15;
				end
				if(in == 4) begin
					state<=5442;
					out<=16;
				end
			end
			3485: begin
				if(in == 0) begin
					state<=3486;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=7375;
					out<=19;
				end
				if(in == 3) begin
					state<=1554;
					out<=20;
				end
				if(in == 4) begin
					state<=5443;
					out<=21;
				end
			end
			3486: begin
				if(in == 0) begin
					state<=3487;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=7376;
					out<=24;
				end
				if(in == 3) begin
					state<=1555;
					out<=25;
				end
				if(in == 4) begin
					state<=5444;
					out<=26;
				end
			end
			3487: begin
				if(in == 0) begin
					state<=3488;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=7377;
					out<=29;
				end
				if(in == 3) begin
					state<=1556;
					out<=30;
				end
				if(in == 4) begin
					state<=5445;
					out<=31;
				end
			end
			3488: begin
				if(in == 0) begin
					state<=3489;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=7378;
					out<=34;
				end
				if(in == 3) begin
					state<=1557;
					out<=35;
				end
				if(in == 4) begin
					state<=5446;
					out<=36;
				end
			end
			3489: begin
				if(in == 0) begin
					state<=3490;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=7379;
					out<=39;
				end
				if(in == 3) begin
					state<=1558;
					out<=40;
				end
				if(in == 4) begin
					state<=5447;
					out<=41;
				end
			end
			3490: begin
				if(in == 0) begin
					state<=3491;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=7380;
					out<=44;
				end
				if(in == 3) begin
					state<=1559;
					out<=45;
				end
				if(in == 4) begin
					state<=5448;
					out<=46;
				end
			end
			3491: begin
				if(in == 0) begin
					state<=3492;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=7381;
					out<=49;
				end
				if(in == 3) begin
					state<=1560;
					out<=50;
				end
				if(in == 4) begin
					state<=5449;
					out<=51;
				end
			end
			3492: begin
				if(in == 0) begin
					state<=3493;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=7382;
					out<=54;
				end
				if(in == 3) begin
					state<=1561;
					out<=55;
				end
				if(in == 4) begin
					state<=5450;
					out<=56;
				end
			end
			3493: begin
				if(in == 0) begin
					state<=3494;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=7383;
					out<=59;
				end
				if(in == 3) begin
					state<=1562;
					out<=60;
				end
				if(in == 4) begin
					state<=5451;
					out<=61;
				end
			end
			3494: begin
				if(in == 0) begin
					state<=3495;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=7384;
					out<=64;
				end
				if(in == 3) begin
					state<=1563;
					out<=65;
				end
				if(in == 4) begin
					state<=5452;
					out<=66;
				end
			end
			3495: begin
				if(in == 0) begin
					state<=3496;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=7385;
					out<=69;
				end
				if(in == 3) begin
					state<=1564;
					out<=70;
				end
				if(in == 4) begin
					state<=5453;
					out<=71;
				end
			end
			3496: begin
				if(in == 0) begin
					state<=3497;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=7386;
					out<=74;
				end
				if(in == 3) begin
					state<=1565;
					out<=75;
				end
				if(in == 4) begin
					state<=5454;
					out<=76;
				end
			end
			3497: begin
				if(in == 0) begin
					state<=3498;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=7387;
					out<=79;
				end
				if(in == 3) begin
					state<=1566;
					out<=80;
				end
				if(in == 4) begin
					state<=5455;
					out<=81;
				end
			end
			3498: begin
				if(in == 0) begin
					state<=3499;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=7388;
					out<=84;
				end
				if(in == 3) begin
					state<=1567;
					out<=85;
				end
				if(in == 4) begin
					state<=5456;
					out<=86;
				end
			end
			3499: begin
				if(in == 0) begin
					state<=3500;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=7389;
					out<=89;
				end
				if(in == 3) begin
					state<=1568;
					out<=90;
				end
				if(in == 4) begin
					state<=5457;
					out<=91;
				end
			end
			3500: begin
				if(in == 0) begin
					state<=3501;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=7390;
					out<=94;
				end
				if(in == 3) begin
					state<=1569;
					out<=95;
				end
				if(in == 4) begin
					state<=5458;
					out<=96;
				end
			end
			3501: begin
				if(in == 0) begin
					state<=3502;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=7391;
					out<=99;
				end
				if(in == 3) begin
					state<=1570;
					out<=100;
				end
				if(in == 4) begin
					state<=5459;
					out<=101;
				end
			end
			3502: begin
				if(in == 0) begin
					state<=3503;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=7392;
					out<=104;
				end
				if(in == 3) begin
					state<=1571;
					out<=105;
				end
				if(in == 4) begin
					state<=5460;
					out<=106;
				end
			end
			3503: begin
				if(in == 0) begin
					state<=3504;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=7393;
					out<=109;
				end
				if(in == 3) begin
					state<=1572;
					out<=110;
				end
				if(in == 4) begin
					state<=5461;
					out<=111;
				end
			end
			3504: begin
				if(in == 0) begin
					state<=3505;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=7394;
					out<=114;
				end
				if(in == 3) begin
					state<=1573;
					out<=115;
				end
				if(in == 4) begin
					state<=5462;
					out<=116;
				end
			end
			3505: begin
				if(in == 0) begin
					state<=3506;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=7395;
					out<=119;
				end
				if(in == 3) begin
					state<=1574;
					out<=120;
				end
				if(in == 4) begin
					state<=5463;
					out<=121;
				end
			end
			3506: begin
				if(in == 0) begin
					state<=3507;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=7396;
					out<=124;
				end
				if(in == 3) begin
					state<=1575;
					out<=125;
				end
				if(in == 4) begin
					state<=5464;
					out<=126;
				end
			end
			3507: begin
				if(in == 0) begin
					state<=3508;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=7397;
					out<=129;
				end
				if(in == 3) begin
					state<=1576;
					out<=130;
				end
				if(in == 4) begin
					state<=5465;
					out<=131;
				end
			end
			3508: begin
				if(in == 0) begin
					state<=2601;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=6490;
					out<=134;
				end
				if(in == 3) begin
					state<=603;
					out<=135;
				end
				if(in == 4) begin
					state<=4501;
					out<=136;
				end
			end
			3509: begin
				if(in == 0) begin
					state<=3510;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=7399;
					out<=139;
				end
				if(in == 3) begin
					state<=1609;
					out<=140;
				end
				if(in == 4) begin
					state<=5498;
					out<=141;
				end
			end
			3510: begin
				if(in == 0) begin
					state<=3511;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=7400;
					out<=144;
				end
				if(in == 3) begin
					state<=1610;
					out<=145;
				end
				if(in == 4) begin
					state<=5499;
					out<=146;
				end
			end
			3511: begin
				if(in == 0) begin
					state<=3512;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=7401;
					out<=149;
				end
				if(in == 3) begin
					state<=1611;
					out<=150;
				end
				if(in == 4) begin
					state<=5500;
					out<=151;
				end
			end
			3512: begin
				if(in == 0) begin
					state<=3513;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=7402;
					out<=154;
				end
				if(in == 3) begin
					state<=1612;
					out<=155;
				end
				if(in == 4) begin
					state<=5501;
					out<=156;
				end
			end
			3513: begin
				if(in == 0) begin
					state<=3514;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=7403;
					out<=159;
				end
				if(in == 3) begin
					state<=1613;
					out<=160;
				end
				if(in == 4) begin
					state<=5502;
					out<=161;
				end
			end
			3514: begin
				if(in == 0) begin
					state<=3515;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=7404;
					out<=164;
				end
				if(in == 3) begin
					state<=1614;
					out<=165;
				end
				if(in == 4) begin
					state<=5503;
					out<=166;
				end
			end
			3515: begin
				if(in == 0) begin
					state<=3516;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=7405;
					out<=169;
				end
				if(in == 3) begin
					state<=1615;
					out<=170;
				end
				if(in == 4) begin
					state<=5504;
					out<=171;
				end
			end
			3516: begin
				if(in == 0) begin
					state<=3517;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=7406;
					out<=174;
				end
				if(in == 3) begin
					state<=1616;
					out<=175;
				end
				if(in == 4) begin
					state<=5505;
					out<=176;
				end
			end
			3517: begin
				if(in == 0) begin
					state<=3518;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=7407;
					out<=179;
				end
				if(in == 3) begin
					state<=1617;
					out<=180;
				end
				if(in == 4) begin
					state<=5506;
					out<=181;
				end
			end
			3518: begin
				if(in == 0) begin
					state<=3519;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=7408;
					out<=184;
				end
				if(in == 3) begin
					state<=1618;
					out<=185;
				end
				if(in == 4) begin
					state<=5507;
					out<=186;
				end
			end
			3519: begin
				if(in == 0) begin
					state<=3520;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=7409;
					out<=189;
				end
				if(in == 3) begin
					state<=1619;
					out<=190;
				end
				if(in == 4) begin
					state<=5508;
					out<=191;
				end
			end
			3520: begin
				if(in == 0) begin
					state<=3521;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=7410;
					out<=194;
				end
				if(in == 3) begin
					state<=1620;
					out<=195;
				end
				if(in == 4) begin
					state<=5509;
					out<=196;
				end
			end
			3521: begin
				if(in == 0) begin
					state<=3522;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=7411;
					out<=199;
				end
				if(in == 3) begin
					state<=1621;
					out<=200;
				end
				if(in == 4) begin
					state<=5510;
					out<=201;
				end
			end
			3522: begin
				if(in == 0) begin
					state<=3523;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=7412;
					out<=204;
				end
				if(in == 3) begin
					state<=1622;
					out<=205;
				end
				if(in == 4) begin
					state<=5511;
					out<=206;
				end
			end
			3523: begin
				if(in == 0) begin
					state<=3524;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=7413;
					out<=209;
				end
				if(in == 3) begin
					state<=1623;
					out<=210;
				end
				if(in == 4) begin
					state<=5512;
					out<=211;
				end
			end
			3524: begin
				if(in == 0) begin
					state<=3525;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=7414;
					out<=214;
				end
				if(in == 3) begin
					state<=1624;
					out<=215;
				end
				if(in == 4) begin
					state<=5513;
					out<=216;
				end
			end
			3525: begin
				if(in == 0) begin
					state<=3526;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=7415;
					out<=219;
				end
				if(in == 3) begin
					state<=1625;
					out<=220;
				end
				if(in == 4) begin
					state<=5514;
					out<=221;
				end
			end
			3526: begin
				if(in == 0) begin
					state<=3527;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=7416;
					out<=224;
				end
				if(in == 3) begin
					state<=1626;
					out<=225;
				end
				if(in == 4) begin
					state<=5515;
					out<=226;
				end
			end
			3527: begin
				if(in == 0) begin
					state<=3528;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=7417;
					out<=229;
				end
				if(in == 3) begin
					state<=1627;
					out<=230;
				end
				if(in == 4) begin
					state<=5516;
					out<=231;
				end
			end
			3528: begin
				if(in == 0) begin
					state<=3529;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=7418;
					out<=234;
				end
				if(in == 3) begin
					state<=1628;
					out<=235;
				end
				if(in == 4) begin
					state<=5517;
					out<=236;
				end
			end
			3529: begin
				if(in == 0) begin
					state<=3530;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=7419;
					out<=239;
				end
				if(in == 3) begin
					state<=1629;
					out<=240;
				end
				if(in == 4) begin
					state<=5518;
					out<=241;
				end
			end
			3530: begin
				if(in == 0) begin
					state<=3531;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=7420;
					out<=244;
				end
				if(in == 3) begin
					state<=1630;
					out<=245;
				end
				if(in == 4) begin
					state<=5519;
					out<=246;
				end
			end
			3531: begin
				if(in == 0) begin
					state<=3532;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=7421;
					out<=249;
				end
				if(in == 3) begin
					state<=1631;
					out<=250;
				end
				if(in == 4) begin
					state<=5520;
					out<=251;
				end
			end
			3532: begin
				if(in == 0) begin
					state<=3533;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=7422;
					out<=254;
				end
				if(in == 3) begin
					state<=1632;
					out<=255;
				end
				if(in == 4) begin
					state<=5521;
					out<=0;
				end
			end
			3533: begin
				if(in == 0) begin
					state<=3534;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=7423;
					out<=3;
				end
				if(in == 3) begin
					state<=1633;
					out<=4;
				end
				if(in == 4) begin
					state<=5522;
					out<=5;
				end
			end
			3534: begin
				if(in == 0) begin
					state<=3535;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=7424;
					out<=8;
				end
				if(in == 3) begin
					state<=1634;
					out<=9;
				end
				if(in == 4) begin
					state<=5523;
					out<=10;
				end
			end
			3535: begin
				if(in == 0) begin
					state<=3536;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=7425;
					out<=13;
				end
				if(in == 3) begin
					state<=1635;
					out<=14;
				end
				if(in == 4) begin
					state<=5524;
					out<=15;
				end
			end
			3536: begin
				if(in == 0) begin
					state<=3537;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=7426;
					out<=18;
				end
				if(in == 3) begin
					state<=1636;
					out<=19;
				end
				if(in == 4) begin
					state<=5525;
					out<=20;
				end
			end
			3537: begin
				if(in == 0) begin
					state<=3538;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=7427;
					out<=23;
				end
				if(in == 3) begin
					state<=1637;
					out<=24;
				end
				if(in == 4) begin
					state<=5526;
					out<=25;
				end
			end
			3538: begin
				if(in == 0) begin
					state<=3539;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=7428;
					out<=28;
				end
				if(in == 3) begin
					state<=1638;
					out<=29;
				end
				if(in == 4) begin
					state<=5527;
					out<=30;
				end
			end
			3539: begin
				if(in == 0) begin
					state<=3540;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=7429;
					out<=33;
				end
				if(in == 3) begin
					state<=1639;
					out<=34;
				end
				if(in == 4) begin
					state<=5528;
					out<=35;
				end
			end
			3540: begin
				if(in == 0) begin
					state<=3541;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=7430;
					out<=38;
				end
				if(in == 3) begin
					state<=1640;
					out<=39;
				end
				if(in == 4) begin
					state<=5529;
					out<=40;
				end
			end
			3541: begin
				if(in == 0) begin
					state<=3542;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=7431;
					out<=43;
				end
				if(in == 3) begin
					state<=1641;
					out<=44;
				end
				if(in == 4) begin
					state<=5530;
					out<=45;
				end
			end
			3542: begin
				if(in == 0) begin
					state<=3543;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=7432;
					out<=48;
				end
				if(in == 3) begin
					state<=1642;
					out<=49;
				end
				if(in == 4) begin
					state<=5531;
					out<=50;
				end
			end
			3543: begin
				if(in == 0) begin
					state<=3544;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=7433;
					out<=53;
				end
				if(in == 3) begin
					state<=1643;
					out<=54;
				end
				if(in == 4) begin
					state<=5532;
					out<=55;
				end
			end
			3544: begin
				if(in == 0) begin
					state<=3545;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=7434;
					out<=58;
				end
				if(in == 3) begin
					state<=1644;
					out<=59;
				end
				if(in == 4) begin
					state<=5533;
					out<=60;
				end
			end
			3545: begin
				if(in == 0) begin
					state<=3546;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=7435;
					out<=63;
				end
				if(in == 3) begin
					state<=1645;
					out<=64;
				end
				if(in == 4) begin
					state<=5534;
					out<=65;
				end
			end
			3546: begin
				if(in == 0) begin
					state<=3547;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=7436;
					out<=68;
				end
				if(in == 3) begin
					state<=1646;
					out<=69;
				end
				if(in == 4) begin
					state<=5535;
					out<=70;
				end
			end
			3547: begin
				if(in == 0) begin
					state<=3548;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=7437;
					out<=73;
				end
				if(in == 3) begin
					state<=1647;
					out<=74;
				end
				if(in == 4) begin
					state<=5536;
					out<=75;
				end
			end
			3548: begin
				if(in == 0) begin
					state<=3549;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=7438;
					out<=78;
				end
				if(in == 3) begin
					state<=1648;
					out<=79;
				end
				if(in == 4) begin
					state<=5537;
					out<=80;
				end
			end
			3549: begin
				if(in == 0) begin
					state<=3550;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=7439;
					out<=83;
				end
				if(in == 3) begin
					state<=1649;
					out<=84;
				end
				if(in == 4) begin
					state<=5538;
					out<=85;
				end
			end
			3550: begin
				if(in == 0) begin
					state<=3551;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=7440;
					out<=88;
				end
				if(in == 3) begin
					state<=1650;
					out<=89;
				end
				if(in == 4) begin
					state<=5539;
					out<=90;
				end
			end
			3551: begin
				if(in == 0) begin
					state<=3552;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=7441;
					out<=93;
				end
				if(in == 3) begin
					state<=1651;
					out<=94;
				end
				if(in == 4) begin
					state<=5540;
					out<=95;
				end
			end
			3552: begin
				if(in == 0) begin
					state<=3553;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=7442;
					out<=98;
				end
				if(in == 3) begin
					state<=1652;
					out<=99;
				end
				if(in == 4) begin
					state<=5541;
					out<=100;
				end
			end
			3553: begin
				if(in == 0) begin
					state<=3554;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=7443;
					out<=103;
				end
				if(in == 3) begin
					state<=1653;
					out<=104;
				end
				if(in == 4) begin
					state<=5542;
					out<=105;
				end
			end
			3554: begin
				if(in == 0) begin
					state<=3555;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=7444;
					out<=108;
				end
				if(in == 3) begin
					state<=1654;
					out<=109;
				end
				if(in == 4) begin
					state<=5543;
					out<=110;
				end
			end
			3555: begin
				if(in == 0) begin
					state<=3556;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=7445;
					out<=113;
				end
				if(in == 3) begin
					state<=1655;
					out<=114;
				end
				if(in == 4) begin
					state<=5544;
					out<=115;
				end
			end
			3556: begin
				if(in == 0) begin
					state<=3557;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=7446;
					out<=118;
				end
				if(in == 3) begin
					state<=1656;
					out<=119;
				end
				if(in == 4) begin
					state<=5545;
					out<=120;
				end
			end
			3557: begin
				if(in == 0) begin
					state<=3558;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=7447;
					out<=123;
				end
				if(in == 3) begin
					state<=1657;
					out<=124;
				end
				if(in == 4) begin
					state<=5546;
					out<=125;
				end
			end
			3558: begin
				if(in == 0) begin
					state<=3559;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=7448;
					out<=128;
				end
				if(in == 3) begin
					state<=1658;
					out<=129;
				end
				if(in == 4) begin
					state<=5547;
					out<=130;
				end
			end
			3559: begin
				if(in == 0) begin
					state<=3560;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=7449;
					out<=133;
				end
				if(in == 3) begin
					state<=1659;
					out<=134;
				end
				if(in == 4) begin
					state<=5548;
					out<=135;
				end
			end
			3560: begin
				if(in == 0) begin
					state<=3561;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=7450;
					out<=138;
				end
				if(in == 3) begin
					state<=1660;
					out<=139;
				end
				if(in == 4) begin
					state<=5549;
					out<=140;
				end
			end
			3561: begin
				if(in == 0) begin
					state<=3562;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=7451;
					out<=143;
				end
				if(in == 3) begin
					state<=1661;
					out<=144;
				end
				if(in == 4) begin
					state<=5550;
					out<=145;
				end
			end
			3562: begin
				if(in == 0) begin
					state<=3563;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=7452;
					out<=148;
				end
				if(in == 3) begin
					state<=1662;
					out<=149;
				end
				if(in == 4) begin
					state<=5551;
					out<=150;
				end
			end
			3563: begin
				if(in == 0) begin
					state<=3564;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=7453;
					out<=153;
				end
				if(in == 3) begin
					state<=1663;
					out<=154;
				end
				if(in == 4) begin
					state<=5552;
					out<=155;
				end
			end
			3564: begin
				if(in == 0) begin
					state<=3565;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=7454;
					out<=158;
				end
				if(in == 3) begin
					state<=1664;
					out<=159;
				end
				if(in == 4) begin
					state<=5553;
					out<=160;
				end
			end
			3565: begin
				if(in == 0) begin
					state<=3566;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=7455;
					out<=163;
				end
				if(in == 3) begin
					state<=1665;
					out<=164;
				end
				if(in == 4) begin
					state<=5554;
					out<=165;
				end
			end
			3566: begin
				if(in == 0) begin
					state<=3567;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=7456;
					out<=168;
				end
				if(in == 3) begin
					state<=1666;
					out<=169;
				end
				if(in == 4) begin
					state<=5555;
					out<=170;
				end
			end
			3567: begin
				if(in == 0) begin
					state<=3568;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=7457;
					out<=173;
				end
				if(in == 3) begin
					state<=1667;
					out<=174;
				end
				if(in == 4) begin
					state<=5556;
					out<=175;
				end
			end
			3568: begin
				if(in == 0) begin
					state<=3569;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=7458;
					out<=178;
				end
				if(in == 3) begin
					state<=1668;
					out<=179;
				end
				if(in == 4) begin
					state<=5557;
					out<=180;
				end
			end
			3569: begin
				if(in == 0) begin
					state<=3570;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=7459;
					out<=183;
				end
				if(in == 3) begin
					state<=1669;
					out<=184;
				end
				if(in == 4) begin
					state<=5558;
					out<=185;
				end
			end
			3570: begin
				if(in == 0) begin
					state<=3571;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=7460;
					out<=188;
				end
				if(in == 3) begin
					state<=1670;
					out<=189;
				end
				if(in == 4) begin
					state<=5559;
					out<=190;
				end
			end
			3571: begin
				if(in == 0) begin
					state<=3572;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=7461;
					out<=193;
				end
				if(in == 3) begin
					state<=1671;
					out<=194;
				end
				if(in == 4) begin
					state<=5560;
					out<=195;
				end
			end
			3572: begin
				if(in == 0) begin
					state<=3573;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=7462;
					out<=198;
				end
				if(in == 3) begin
					state<=1672;
					out<=199;
				end
				if(in == 4) begin
					state<=5561;
					out<=200;
				end
			end
			3573: begin
				if(in == 0) begin
					state<=3574;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=7463;
					out<=203;
				end
				if(in == 3) begin
					state<=1673;
					out<=204;
				end
				if(in == 4) begin
					state<=5562;
					out<=205;
				end
			end
			3574: begin
				if(in == 0) begin
					state<=3575;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=7464;
					out<=208;
				end
				if(in == 3) begin
					state<=1674;
					out<=209;
				end
				if(in == 4) begin
					state<=5563;
					out<=210;
				end
			end
			3575: begin
				if(in == 0) begin
					state<=3576;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=7465;
					out<=213;
				end
				if(in == 3) begin
					state<=1675;
					out<=214;
				end
				if(in == 4) begin
					state<=5564;
					out<=215;
				end
			end
			3576: begin
				if(in == 0) begin
					state<=3577;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=7466;
					out<=218;
				end
				if(in == 3) begin
					state<=1676;
					out<=219;
				end
				if(in == 4) begin
					state<=5565;
					out<=220;
				end
			end
			3577: begin
				if(in == 0) begin
					state<=3578;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=7467;
					out<=223;
				end
				if(in == 3) begin
					state<=1677;
					out<=224;
				end
				if(in == 4) begin
					state<=5566;
					out<=225;
				end
			end
			3578: begin
				if(in == 0) begin
					state<=3579;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=7468;
					out<=228;
				end
				if(in == 3) begin
					state<=1678;
					out<=229;
				end
				if(in == 4) begin
					state<=5567;
					out<=230;
				end
			end
			3579: begin
				if(in == 0) begin
					state<=3580;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=7469;
					out<=233;
				end
				if(in == 3) begin
					state<=1679;
					out<=234;
				end
				if(in == 4) begin
					state<=5568;
					out<=235;
				end
			end
			3580: begin
				if(in == 0) begin
					state<=3581;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=7470;
					out<=238;
				end
				if(in == 3) begin
					state<=1680;
					out<=239;
				end
				if(in == 4) begin
					state<=5569;
					out<=240;
				end
			end
			3581: begin
				if(in == 0) begin
					state<=3582;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=7471;
					out<=243;
				end
				if(in == 3) begin
					state<=1681;
					out<=244;
				end
				if(in == 4) begin
					state<=5570;
					out<=245;
				end
			end
			3582: begin
				if(in == 0) begin
					state<=3583;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=7472;
					out<=248;
				end
				if(in == 3) begin
					state<=1682;
					out<=249;
				end
				if(in == 4) begin
					state<=5571;
					out<=250;
				end
			end
			3583: begin
				if(in == 0) begin
					state<=3584;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=7473;
					out<=253;
				end
				if(in == 3) begin
					state<=1683;
					out<=254;
				end
				if(in == 4) begin
					state<=5572;
					out<=255;
				end
			end
			3584: begin
				if(in == 0) begin
					state<=3585;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=7474;
					out<=2;
				end
				if(in == 3) begin
					state<=1684;
					out<=3;
				end
				if(in == 4) begin
					state<=5573;
					out<=4;
				end
			end
			3585: begin
				if(in == 0) begin
					state<=3586;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=7475;
					out<=7;
				end
				if(in == 3) begin
					state<=1685;
					out<=8;
				end
				if(in == 4) begin
					state<=5574;
					out<=9;
				end
			end
			3586: begin
				if(in == 0) begin
					state<=3587;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=7476;
					out<=12;
				end
				if(in == 3) begin
					state<=1686;
					out<=13;
				end
				if(in == 4) begin
					state<=5575;
					out<=14;
				end
			end
			3587: begin
				if(in == 0) begin
					state<=3588;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=7477;
					out<=17;
				end
				if(in == 3) begin
					state<=1687;
					out<=18;
				end
				if(in == 4) begin
					state<=5576;
					out<=19;
				end
			end
			3588: begin
				if(in == 0) begin
					state<=3589;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=7478;
					out<=22;
				end
				if(in == 3) begin
					state<=1688;
					out<=23;
				end
				if(in == 4) begin
					state<=5577;
					out<=24;
				end
			end
			3589: begin
				if(in == 0) begin
					state<=3590;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=7479;
					out<=27;
				end
				if(in == 3) begin
					state<=1689;
					out<=28;
				end
				if(in == 4) begin
					state<=5578;
					out<=29;
				end
			end
			3590: begin
				if(in == 0) begin
					state<=3591;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=7480;
					out<=32;
				end
				if(in == 3) begin
					state<=1690;
					out<=33;
				end
				if(in == 4) begin
					state<=5579;
					out<=34;
				end
			end
			3591: begin
				if(in == 0) begin
					state<=3592;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=7481;
					out<=37;
				end
				if(in == 3) begin
					state<=1691;
					out<=38;
				end
				if(in == 4) begin
					state<=5580;
					out<=39;
				end
			end
			3592: begin
				if(in == 0) begin
					state<=3593;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=7482;
					out<=42;
				end
				if(in == 3) begin
					state<=1692;
					out<=43;
				end
				if(in == 4) begin
					state<=5581;
					out<=44;
				end
			end
			3593: begin
				if(in == 0) begin
					state<=3594;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=7483;
					out<=47;
				end
				if(in == 3) begin
					state<=1693;
					out<=48;
				end
				if(in == 4) begin
					state<=5582;
					out<=49;
				end
			end
			3594: begin
				if(in == 0) begin
					state<=3595;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=7484;
					out<=52;
				end
				if(in == 3) begin
					state<=1694;
					out<=53;
				end
				if(in == 4) begin
					state<=5583;
					out<=54;
				end
			end
			3595: begin
				if(in == 0) begin
					state<=3596;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=7485;
					out<=57;
				end
				if(in == 3) begin
					state<=1695;
					out<=58;
				end
				if(in == 4) begin
					state<=5584;
					out<=59;
				end
			end
			3596: begin
				if(in == 0) begin
					state<=3597;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=7486;
					out<=62;
				end
				if(in == 3) begin
					state<=1696;
					out<=63;
				end
				if(in == 4) begin
					state<=5585;
					out<=64;
				end
			end
			3597: begin
				if(in == 0) begin
					state<=3598;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=7487;
					out<=67;
				end
				if(in == 3) begin
					state<=1697;
					out<=68;
				end
				if(in == 4) begin
					state<=5586;
					out<=69;
				end
			end
			3598: begin
				if(in == 0) begin
					state<=3599;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=7488;
					out<=72;
				end
				if(in == 3) begin
					state<=1698;
					out<=73;
				end
				if(in == 4) begin
					state<=5587;
					out<=74;
				end
			end
			3599: begin
				if(in == 0) begin
					state<=3600;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=7489;
					out<=77;
				end
				if(in == 3) begin
					state<=1699;
					out<=78;
				end
				if(in == 4) begin
					state<=5588;
					out<=79;
				end
			end
			3600: begin
				if(in == 0) begin
					state<=3601;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=7490;
					out<=82;
				end
				if(in == 3) begin
					state<=1700;
					out<=83;
				end
				if(in == 4) begin
					state<=5589;
					out<=84;
				end
			end
			3601: begin
				if(in == 0) begin
					state<=3602;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=7491;
					out<=87;
				end
				if(in == 3) begin
					state<=1701;
					out<=88;
				end
				if(in == 4) begin
					state<=5590;
					out<=89;
				end
			end
			3602: begin
				if(in == 0) begin
					state<=3603;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=7492;
					out<=92;
				end
				if(in == 3) begin
					state<=1702;
					out<=93;
				end
				if(in == 4) begin
					state<=5591;
					out<=94;
				end
			end
			3603: begin
				if(in == 0) begin
					state<=3604;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=7493;
					out<=97;
				end
				if(in == 3) begin
					state<=1703;
					out<=98;
				end
				if(in == 4) begin
					state<=5592;
					out<=99;
				end
			end
			3604: begin
				if(in == 0) begin
					state<=3605;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=7494;
					out<=102;
				end
				if(in == 3) begin
					state<=1704;
					out<=103;
				end
				if(in == 4) begin
					state<=5593;
					out<=104;
				end
			end
			3605: begin
				if(in == 0) begin
					state<=3606;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=7495;
					out<=107;
				end
				if(in == 3) begin
					state<=1705;
					out<=108;
				end
				if(in == 4) begin
					state<=5594;
					out<=109;
				end
			end
			3606: begin
				if(in == 0) begin
					state<=3607;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=7496;
					out<=112;
				end
				if(in == 3) begin
					state<=1706;
					out<=113;
				end
				if(in == 4) begin
					state<=5595;
					out<=114;
				end
			end
			3607: begin
				if(in == 0) begin
					state<=3608;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=7497;
					out<=117;
				end
				if(in == 3) begin
					state<=1707;
					out<=118;
				end
				if(in == 4) begin
					state<=5596;
					out<=119;
				end
			end
			3608: begin
				if(in == 0) begin
					state<=3609;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=7498;
					out<=122;
				end
				if(in == 3) begin
					state<=1708;
					out<=123;
				end
				if(in == 4) begin
					state<=5597;
					out<=124;
				end
			end
			3609: begin
				if(in == 0) begin
					state<=3610;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=7499;
					out<=127;
				end
				if(in == 3) begin
					state<=1709;
					out<=128;
				end
				if(in == 4) begin
					state<=5598;
					out<=129;
				end
			end
			3610: begin
				if(in == 0) begin
					state<=3611;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=7500;
					out<=132;
				end
				if(in == 3) begin
					state<=1710;
					out<=133;
				end
				if(in == 4) begin
					state<=5599;
					out<=134;
				end
			end
			3611: begin
				if(in == 0) begin
					state<=3612;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=7501;
					out<=137;
				end
				if(in == 3) begin
					state<=1711;
					out<=138;
				end
				if(in == 4) begin
					state<=5600;
					out<=139;
				end
			end
			3612: begin
				if(in == 0) begin
					state<=3613;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=7502;
					out<=142;
				end
				if(in == 3) begin
					state<=1712;
					out<=143;
				end
				if(in == 4) begin
					state<=5601;
					out<=144;
				end
			end
			3613: begin
				if(in == 0) begin
					state<=3614;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=7503;
					out<=147;
				end
				if(in == 3) begin
					state<=1713;
					out<=148;
				end
				if(in == 4) begin
					state<=5602;
					out<=149;
				end
			end
			3614: begin
				if(in == 0) begin
					state<=3615;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=7504;
					out<=152;
				end
				if(in == 3) begin
					state<=1714;
					out<=153;
				end
				if(in == 4) begin
					state<=5603;
					out<=154;
				end
			end
			3615: begin
				if(in == 0) begin
					state<=3616;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=7505;
					out<=157;
				end
				if(in == 3) begin
					state<=1715;
					out<=158;
				end
				if(in == 4) begin
					state<=5604;
					out<=159;
				end
			end
			3616: begin
				if(in == 0) begin
					state<=3617;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=7506;
					out<=162;
				end
				if(in == 3) begin
					state<=1716;
					out<=163;
				end
				if(in == 4) begin
					state<=5605;
					out<=164;
				end
			end
			3617: begin
				if(in == 0) begin
					state<=3618;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=7507;
					out<=167;
				end
				if(in == 3) begin
					state<=1717;
					out<=168;
				end
				if(in == 4) begin
					state<=5606;
					out<=169;
				end
			end
			3618: begin
				if(in == 0) begin
					state<=3619;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=7508;
					out<=172;
				end
				if(in == 3) begin
					state<=1718;
					out<=173;
				end
				if(in == 4) begin
					state<=5607;
					out<=174;
				end
			end
			3619: begin
				if(in == 0) begin
					state<=3620;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=7509;
					out<=177;
				end
				if(in == 3) begin
					state<=1719;
					out<=178;
				end
				if(in == 4) begin
					state<=5608;
					out<=179;
				end
			end
			3620: begin
				if(in == 0) begin
					state<=3621;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=7510;
					out<=182;
				end
				if(in == 3) begin
					state<=1720;
					out<=183;
				end
				if(in == 4) begin
					state<=5609;
					out<=184;
				end
			end
			3621: begin
				if(in == 0) begin
					state<=3622;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=7511;
					out<=187;
				end
				if(in == 3) begin
					state<=1721;
					out<=188;
				end
				if(in == 4) begin
					state<=5610;
					out<=189;
				end
			end
			3622: begin
				if(in == 0) begin
					state<=3623;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=7512;
					out<=192;
				end
				if(in == 3) begin
					state<=1722;
					out<=193;
				end
				if(in == 4) begin
					state<=5611;
					out<=194;
				end
			end
			3623: begin
				if(in == 0) begin
					state<=3624;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=7513;
					out<=197;
				end
				if(in == 3) begin
					state<=1723;
					out<=198;
				end
				if(in == 4) begin
					state<=5612;
					out<=199;
				end
			end
			3624: begin
				if(in == 0) begin
					state<=3625;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=7514;
					out<=202;
				end
				if(in == 3) begin
					state<=1724;
					out<=203;
				end
				if(in == 4) begin
					state<=5613;
					out<=204;
				end
			end
			3625: begin
				if(in == 0) begin
					state<=3626;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=7515;
					out<=207;
				end
				if(in == 3) begin
					state<=1725;
					out<=208;
				end
				if(in == 4) begin
					state<=5614;
					out<=209;
				end
			end
			3626: begin
				if(in == 0) begin
					state<=3627;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=7516;
					out<=212;
				end
				if(in == 3) begin
					state<=1726;
					out<=213;
				end
				if(in == 4) begin
					state<=5615;
					out<=214;
				end
			end
			3627: begin
				if(in == 0) begin
					state<=3628;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=7517;
					out<=217;
				end
				if(in == 3) begin
					state<=1727;
					out<=218;
				end
				if(in == 4) begin
					state<=5616;
					out<=219;
				end
			end
			3628: begin
				if(in == 0) begin
					state<=3629;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=7518;
					out<=222;
				end
				if(in == 3) begin
					state<=1728;
					out<=223;
				end
				if(in == 4) begin
					state<=5617;
					out<=224;
				end
			end
			3629: begin
				if(in == 0) begin
					state<=3630;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=7519;
					out<=227;
				end
				if(in == 3) begin
					state<=1729;
					out<=228;
				end
				if(in == 4) begin
					state<=5618;
					out<=229;
				end
			end
			3630: begin
				if(in == 0) begin
					state<=3631;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=7520;
					out<=232;
				end
				if(in == 3) begin
					state<=1730;
					out<=233;
				end
				if(in == 4) begin
					state<=5619;
					out<=234;
				end
			end
			3631: begin
				if(in == 0) begin
					state<=3632;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=7521;
					out<=237;
				end
				if(in == 3) begin
					state<=1731;
					out<=238;
				end
				if(in == 4) begin
					state<=5620;
					out<=239;
				end
			end
			3632: begin
				if(in == 0) begin
					state<=3633;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=7522;
					out<=242;
				end
				if(in == 3) begin
					state<=1732;
					out<=243;
				end
				if(in == 4) begin
					state<=5621;
					out<=244;
				end
			end
			3633: begin
				if(in == 0) begin
					state<=3634;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=7523;
					out<=247;
				end
				if(in == 3) begin
					state<=1733;
					out<=248;
				end
				if(in == 4) begin
					state<=5622;
					out<=249;
				end
			end
			3634: begin
				if(in == 0) begin
					state<=3635;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=7524;
					out<=252;
				end
				if(in == 3) begin
					state<=1734;
					out<=253;
				end
				if(in == 4) begin
					state<=5623;
					out<=254;
				end
			end
			3635: begin
				if(in == 0) begin
					state<=3636;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=7525;
					out<=1;
				end
				if(in == 3) begin
					state<=1735;
					out<=2;
				end
				if(in == 4) begin
					state<=5624;
					out<=3;
				end
			end
			3636: begin
				if(in == 0) begin
					state<=3637;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=7526;
					out<=6;
				end
				if(in == 3) begin
					state<=1736;
					out<=7;
				end
				if(in == 4) begin
					state<=5625;
					out<=8;
				end
			end
			3637: begin
				if(in == 0) begin
					state<=3638;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=7527;
					out<=11;
				end
				if(in == 3) begin
					state<=1737;
					out<=12;
				end
				if(in == 4) begin
					state<=5626;
					out<=13;
				end
			end
			3638: begin
				if(in == 0) begin
					state<=3639;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=7528;
					out<=16;
				end
				if(in == 3) begin
					state<=1738;
					out<=17;
				end
				if(in == 4) begin
					state<=5627;
					out<=18;
				end
			end
			3639: begin
				if(in == 0) begin
					state<=3640;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=7529;
					out<=21;
				end
				if(in == 3) begin
					state<=1739;
					out<=22;
				end
				if(in == 4) begin
					state<=5628;
					out<=23;
				end
			end
			3640: begin
				if(in == 0) begin
					state<=3641;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=7530;
					out<=26;
				end
				if(in == 3) begin
					state<=1740;
					out<=27;
				end
				if(in == 4) begin
					state<=5629;
					out<=28;
				end
			end
			3641: begin
				if(in == 0) begin
					state<=3642;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=7531;
					out<=31;
				end
				if(in == 3) begin
					state<=1741;
					out<=32;
				end
				if(in == 4) begin
					state<=5630;
					out<=33;
				end
			end
			3642: begin
				if(in == 0) begin
					state<=3643;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=7532;
					out<=36;
				end
				if(in == 3) begin
					state<=1742;
					out<=37;
				end
				if(in == 4) begin
					state<=5631;
					out<=38;
				end
			end
			3643: begin
				if(in == 0) begin
					state<=3644;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=7533;
					out<=41;
				end
				if(in == 3) begin
					state<=1743;
					out<=42;
				end
				if(in == 4) begin
					state<=5632;
					out<=43;
				end
			end
			3644: begin
				if(in == 0) begin
					state<=3645;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=7534;
					out<=46;
				end
				if(in == 3) begin
					state<=1744;
					out<=47;
				end
				if(in == 4) begin
					state<=5633;
					out<=48;
				end
			end
			3645: begin
				if(in == 0) begin
					state<=3646;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=7535;
					out<=51;
				end
				if(in == 3) begin
					state<=1745;
					out<=52;
				end
				if(in == 4) begin
					state<=5634;
					out<=53;
				end
			end
			3646: begin
				if(in == 0) begin
					state<=3647;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=7536;
					out<=56;
				end
				if(in == 3) begin
					state<=1746;
					out<=57;
				end
				if(in == 4) begin
					state<=5635;
					out<=58;
				end
			end
			3647: begin
				if(in == 0) begin
					state<=3648;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=7537;
					out<=61;
				end
				if(in == 3) begin
					state<=1747;
					out<=62;
				end
				if(in == 4) begin
					state<=5636;
					out<=63;
				end
			end
			3648: begin
				if(in == 0) begin
					state<=3649;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=7538;
					out<=66;
				end
				if(in == 3) begin
					state<=1748;
					out<=67;
				end
				if(in == 4) begin
					state<=5637;
					out<=68;
				end
			end
			3649: begin
				if(in == 0) begin
					state<=3650;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=7539;
					out<=71;
				end
				if(in == 3) begin
					state<=1749;
					out<=72;
				end
				if(in == 4) begin
					state<=5638;
					out<=73;
				end
			end
			3650: begin
				if(in == 0) begin
					state<=3651;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=7540;
					out<=76;
				end
				if(in == 3) begin
					state<=1750;
					out<=77;
				end
				if(in == 4) begin
					state<=5639;
					out<=78;
				end
			end
			3651: begin
				if(in == 0) begin
					state<=3652;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=7541;
					out<=81;
				end
				if(in == 3) begin
					state<=1751;
					out<=82;
				end
				if(in == 4) begin
					state<=5640;
					out<=83;
				end
			end
			3652: begin
				if(in == 0) begin
					state<=3653;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=7542;
					out<=86;
				end
				if(in == 3) begin
					state<=1752;
					out<=87;
				end
				if(in == 4) begin
					state<=5641;
					out<=88;
				end
			end
			3653: begin
				if(in == 0) begin
					state<=3654;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=7543;
					out<=91;
				end
				if(in == 3) begin
					state<=1753;
					out<=92;
				end
				if(in == 4) begin
					state<=5642;
					out<=93;
				end
			end
			3654: begin
				if(in == 0) begin
					state<=3655;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=7544;
					out<=96;
				end
				if(in == 3) begin
					state<=1754;
					out<=97;
				end
				if(in == 4) begin
					state<=5643;
					out<=98;
				end
			end
			3655: begin
				if(in == 0) begin
					state<=3656;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=7545;
					out<=101;
				end
				if(in == 3) begin
					state<=1755;
					out<=102;
				end
				if(in == 4) begin
					state<=5644;
					out<=103;
				end
			end
			3656: begin
				if(in == 0) begin
					state<=3657;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=7546;
					out<=106;
				end
				if(in == 3) begin
					state<=1756;
					out<=107;
				end
				if(in == 4) begin
					state<=5645;
					out<=108;
				end
			end
			3657: begin
				if(in == 0) begin
					state<=3658;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=7547;
					out<=111;
				end
				if(in == 3) begin
					state<=1757;
					out<=112;
				end
				if(in == 4) begin
					state<=5646;
					out<=113;
				end
			end
			3658: begin
				if(in == 0) begin
					state<=3659;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=7548;
					out<=116;
				end
				if(in == 3) begin
					state<=1758;
					out<=117;
				end
				if(in == 4) begin
					state<=5647;
					out<=118;
				end
			end
			3659: begin
				if(in == 0) begin
					state<=3660;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=7549;
					out<=121;
				end
				if(in == 3) begin
					state<=1759;
					out<=122;
				end
				if(in == 4) begin
					state<=5648;
					out<=123;
				end
			end
			3660: begin
				if(in == 0) begin
					state<=3661;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=7550;
					out<=126;
				end
				if(in == 3) begin
					state<=1760;
					out<=127;
				end
				if(in == 4) begin
					state<=5649;
					out<=128;
				end
			end
			3661: begin
				if(in == 0) begin
					state<=3662;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=7551;
					out<=131;
				end
				if(in == 3) begin
					state<=1761;
					out<=132;
				end
				if(in == 4) begin
					state<=5650;
					out<=133;
				end
			end
			3662: begin
				if(in == 0) begin
					state<=3663;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=7552;
					out<=136;
				end
				if(in == 3) begin
					state<=1762;
					out<=137;
				end
				if(in == 4) begin
					state<=5651;
					out<=138;
				end
			end
			3663: begin
				if(in == 0) begin
					state<=3664;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=7553;
					out<=141;
				end
				if(in == 3) begin
					state<=1763;
					out<=142;
				end
				if(in == 4) begin
					state<=5652;
					out<=143;
				end
			end
			3664: begin
				if(in == 0) begin
					state<=3665;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=7554;
					out<=146;
				end
				if(in == 3) begin
					state<=1764;
					out<=147;
				end
				if(in == 4) begin
					state<=5653;
					out<=148;
				end
			end
			3665: begin
				if(in == 0) begin
					state<=3666;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=7555;
					out<=151;
				end
				if(in == 3) begin
					state<=1765;
					out<=152;
				end
				if(in == 4) begin
					state<=5654;
					out<=153;
				end
			end
			3666: begin
				if(in == 0) begin
					state<=3667;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=7556;
					out<=156;
				end
				if(in == 3) begin
					state<=1766;
					out<=157;
				end
				if(in == 4) begin
					state<=5655;
					out<=158;
				end
			end
			3667: begin
				if(in == 0) begin
					state<=3668;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=7557;
					out<=161;
				end
				if(in == 3) begin
					state<=1767;
					out<=162;
				end
				if(in == 4) begin
					state<=5656;
					out<=163;
				end
			end
			3668: begin
				if(in == 0) begin
					state<=3669;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=7558;
					out<=166;
				end
				if(in == 3) begin
					state<=1768;
					out<=167;
				end
				if(in == 4) begin
					state<=5657;
					out<=168;
				end
			end
			3669: begin
				if(in == 0) begin
					state<=3670;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=7559;
					out<=171;
				end
				if(in == 3) begin
					state<=1769;
					out<=172;
				end
				if(in == 4) begin
					state<=5658;
					out<=173;
				end
			end
			3670: begin
				if(in == 0) begin
					state<=3671;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=7560;
					out<=176;
				end
				if(in == 3) begin
					state<=1770;
					out<=177;
				end
				if(in == 4) begin
					state<=5659;
					out<=178;
				end
			end
			3671: begin
				if(in == 0) begin
					state<=3672;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=7561;
					out<=181;
				end
				if(in == 3) begin
					state<=1771;
					out<=182;
				end
				if(in == 4) begin
					state<=5660;
					out<=183;
				end
			end
			3672: begin
				if(in == 0) begin
					state<=3673;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=7562;
					out<=186;
				end
				if(in == 3) begin
					state<=1772;
					out<=187;
				end
				if(in == 4) begin
					state<=5661;
					out<=188;
				end
			end
			3673: begin
				if(in == 0) begin
					state<=3674;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=7563;
					out<=191;
				end
				if(in == 3) begin
					state<=1773;
					out<=192;
				end
				if(in == 4) begin
					state<=5662;
					out<=193;
				end
			end
			3674: begin
				if(in == 0) begin
					state<=3675;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=7564;
					out<=196;
				end
				if(in == 3) begin
					state<=1774;
					out<=197;
				end
				if(in == 4) begin
					state<=5663;
					out<=198;
				end
			end
			3675: begin
				if(in == 0) begin
					state<=3676;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=7565;
					out<=201;
				end
				if(in == 3) begin
					state<=1775;
					out<=202;
				end
				if(in == 4) begin
					state<=5664;
					out<=203;
				end
			end
			3676: begin
				if(in == 0) begin
					state<=3677;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=7566;
					out<=206;
				end
				if(in == 3) begin
					state<=1776;
					out<=207;
				end
				if(in == 4) begin
					state<=5665;
					out<=208;
				end
			end
			3677: begin
				if(in == 0) begin
					state<=3678;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=7567;
					out<=211;
				end
				if(in == 3) begin
					state<=1777;
					out<=212;
				end
				if(in == 4) begin
					state<=5666;
					out<=213;
				end
			end
			3678: begin
				if(in == 0) begin
					state<=3679;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=7568;
					out<=216;
				end
				if(in == 3) begin
					state<=1778;
					out<=217;
				end
				if(in == 4) begin
					state<=5667;
					out<=218;
				end
			end
			3679: begin
				if(in == 0) begin
					state<=3680;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=7569;
					out<=221;
				end
				if(in == 3) begin
					state<=1779;
					out<=222;
				end
				if(in == 4) begin
					state<=5668;
					out<=223;
				end
			end
			3680: begin
				if(in == 0) begin
					state<=3681;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=7570;
					out<=226;
				end
				if(in == 3) begin
					state<=1780;
					out<=227;
				end
				if(in == 4) begin
					state<=5669;
					out<=228;
				end
			end
			3681: begin
				if(in == 0) begin
					state<=3682;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=7571;
					out<=231;
				end
				if(in == 3) begin
					state<=1781;
					out<=232;
				end
				if(in == 4) begin
					state<=5670;
					out<=233;
				end
			end
			3682: begin
				if(in == 0) begin
					state<=3683;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=7572;
					out<=236;
				end
				if(in == 3) begin
					state<=1782;
					out<=237;
				end
				if(in == 4) begin
					state<=5671;
					out<=238;
				end
			end
			3683: begin
				if(in == 0) begin
					state<=3684;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=7573;
					out<=241;
				end
				if(in == 3) begin
					state<=1783;
					out<=242;
				end
				if(in == 4) begin
					state<=5672;
					out<=243;
				end
			end
			3684: begin
				if(in == 0) begin
					state<=3685;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=7574;
					out<=246;
				end
				if(in == 3) begin
					state<=1784;
					out<=247;
				end
				if(in == 4) begin
					state<=5673;
					out<=248;
				end
			end
			3685: begin
				if(in == 0) begin
					state<=3686;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=7575;
					out<=251;
				end
				if(in == 3) begin
					state<=1785;
					out<=252;
				end
				if(in == 4) begin
					state<=5674;
					out<=253;
				end
			end
			3686: begin
				if(in == 0) begin
					state<=3687;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=7576;
					out<=0;
				end
				if(in == 3) begin
					state<=1786;
					out<=1;
				end
				if(in == 4) begin
					state<=5675;
					out<=2;
				end
			end
			3687: begin
				if(in == 0) begin
					state<=3688;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=7577;
					out<=5;
				end
				if(in == 3) begin
					state<=1787;
					out<=6;
				end
				if(in == 4) begin
					state<=5676;
					out<=7;
				end
			end
			3688: begin
				if(in == 0) begin
					state<=3689;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=7578;
					out<=10;
				end
				if(in == 3) begin
					state<=1788;
					out<=11;
				end
				if(in == 4) begin
					state<=5677;
					out<=12;
				end
			end
			3689: begin
				if(in == 0) begin
					state<=3690;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=7579;
					out<=15;
				end
				if(in == 3) begin
					state<=1789;
					out<=16;
				end
				if(in == 4) begin
					state<=5678;
					out<=17;
				end
			end
			3690: begin
				if(in == 0) begin
					state<=3691;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=7580;
					out<=20;
				end
				if(in == 3) begin
					state<=1790;
					out<=21;
				end
				if(in == 4) begin
					state<=5679;
					out<=22;
				end
			end
			3691: begin
				if(in == 0) begin
					state<=3692;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=7581;
					out<=25;
				end
				if(in == 3) begin
					state<=1791;
					out<=26;
				end
				if(in == 4) begin
					state<=5680;
					out<=27;
				end
			end
			3692: begin
				if(in == 0) begin
					state<=3693;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=7582;
					out<=30;
				end
				if(in == 3) begin
					state<=1792;
					out<=31;
				end
				if(in == 4) begin
					state<=5681;
					out<=32;
				end
			end
			3693: begin
				if(in == 0) begin
					state<=3694;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=7583;
					out<=35;
				end
				if(in == 3) begin
					state<=1793;
					out<=36;
				end
				if(in == 4) begin
					state<=5682;
					out<=37;
				end
			end
			3694: begin
				if(in == 0) begin
					state<=3695;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=7584;
					out<=40;
				end
				if(in == 3) begin
					state<=1794;
					out<=41;
				end
				if(in == 4) begin
					state<=5683;
					out<=42;
				end
			end
			3695: begin
				if(in == 0) begin
					state<=3696;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=7585;
					out<=45;
				end
				if(in == 3) begin
					state<=1795;
					out<=46;
				end
				if(in == 4) begin
					state<=5684;
					out<=47;
				end
			end
			3696: begin
				if(in == 0) begin
					state<=3697;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=7586;
					out<=50;
				end
				if(in == 3) begin
					state<=1796;
					out<=51;
				end
				if(in == 4) begin
					state<=5685;
					out<=52;
				end
			end
			3697: begin
				if(in == 0) begin
					state<=3698;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=7587;
					out<=55;
				end
				if(in == 3) begin
					state<=1797;
					out<=56;
				end
				if(in == 4) begin
					state<=5686;
					out<=57;
				end
			end
			3698: begin
				if(in == 0) begin
					state<=3699;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=7588;
					out<=60;
				end
				if(in == 3) begin
					state<=1798;
					out<=61;
				end
				if(in == 4) begin
					state<=5687;
					out<=62;
				end
			end
			3699: begin
				if(in == 0) begin
					state<=3700;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=7589;
					out<=65;
				end
				if(in == 3) begin
					state<=1799;
					out<=66;
				end
				if(in == 4) begin
					state<=5688;
					out<=67;
				end
			end
			3700: begin
				if(in == 0) begin
					state<=3701;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=7590;
					out<=70;
				end
				if(in == 3) begin
					state<=1800;
					out<=71;
				end
				if(in == 4) begin
					state<=5689;
					out<=72;
				end
			end
			3701: begin
				if(in == 0) begin
					state<=3702;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=7591;
					out<=75;
				end
				if(in == 3) begin
					state<=1801;
					out<=76;
				end
				if(in == 4) begin
					state<=5690;
					out<=77;
				end
			end
			3702: begin
				if(in == 0) begin
					state<=3703;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=7592;
					out<=80;
				end
				if(in == 3) begin
					state<=1802;
					out<=81;
				end
				if(in == 4) begin
					state<=5691;
					out<=82;
				end
			end
			3703: begin
				if(in == 0) begin
					state<=3704;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=7593;
					out<=85;
				end
				if(in == 3) begin
					state<=1803;
					out<=86;
				end
				if(in == 4) begin
					state<=5692;
					out<=87;
				end
			end
			3704: begin
				if(in == 0) begin
					state<=3705;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=7594;
					out<=90;
				end
				if(in == 3) begin
					state<=1804;
					out<=91;
				end
				if(in == 4) begin
					state<=5693;
					out<=92;
				end
			end
			3705: begin
				if(in == 0) begin
					state<=3706;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=7595;
					out<=95;
				end
				if(in == 3) begin
					state<=1805;
					out<=96;
				end
				if(in == 4) begin
					state<=5694;
					out<=97;
				end
			end
			3706: begin
				if(in == 0) begin
					state<=3707;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=7596;
					out<=100;
				end
				if(in == 3) begin
					state<=1806;
					out<=101;
				end
				if(in == 4) begin
					state<=5695;
					out<=102;
				end
			end
			3707: begin
				if(in == 0) begin
					state<=3708;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=7597;
					out<=105;
				end
				if(in == 3) begin
					state<=1807;
					out<=106;
				end
				if(in == 4) begin
					state<=5696;
					out<=107;
				end
			end
			3708: begin
				if(in == 0) begin
					state<=3709;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=7598;
					out<=110;
				end
				if(in == 3) begin
					state<=1808;
					out<=111;
				end
				if(in == 4) begin
					state<=5697;
					out<=112;
				end
			end
			3709: begin
				if(in == 0) begin
					state<=3710;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=7599;
					out<=115;
				end
				if(in == 3) begin
					state<=1809;
					out<=116;
				end
				if(in == 4) begin
					state<=5698;
					out<=117;
				end
			end
			3710: begin
				if(in == 0) begin
					state<=3711;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=7600;
					out<=120;
				end
				if(in == 3) begin
					state<=1810;
					out<=121;
				end
				if(in == 4) begin
					state<=5699;
					out<=122;
				end
			end
			3711: begin
				if(in == 0) begin
					state<=3712;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=7601;
					out<=125;
				end
				if(in == 3) begin
					state<=1811;
					out<=126;
				end
				if(in == 4) begin
					state<=5700;
					out<=127;
				end
			end
			3712: begin
				if(in == 0) begin
					state<=3713;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=7602;
					out<=130;
				end
				if(in == 3) begin
					state<=1812;
					out<=131;
				end
				if(in == 4) begin
					state<=5701;
					out<=132;
				end
			end
			3713: begin
				if(in == 0) begin
					state<=3714;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=7603;
					out<=135;
				end
				if(in == 3) begin
					state<=1813;
					out<=136;
				end
				if(in == 4) begin
					state<=5702;
					out<=137;
				end
			end
			3714: begin
				if(in == 0) begin
					state<=3715;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=7604;
					out<=140;
				end
				if(in == 3) begin
					state<=1814;
					out<=141;
				end
				if(in == 4) begin
					state<=5703;
					out<=142;
				end
			end
			3715: begin
				if(in == 0) begin
					state<=3716;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=7605;
					out<=145;
				end
				if(in == 3) begin
					state<=1815;
					out<=146;
				end
				if(in == 4) begin
					state<=5704;
					out<=147;
				end
			end
			3716: begin
				if(in == 0) begin
					state<=3717;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=7606;
					out<=150;
				end
				if(in == 3) begin
					state<=1816;
					out<=151;
				end
				if(in == 4) begin
					state<=5705;
					out<=152;
				end
			end
			3717: begin
				if(in == 0) begin
					state<=3718;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=7607;
					out<=155;
				end
				if(in == 3) begin
					state<=1817;
					out<=156;
				end
				if(in == 4) begin
					state<=5706;
					out<=157;
				end
			end
			3718: begin
				if(in == 0) begin
					state<=3719;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=7608;
					out<=160;
				end
				if(in == 3) begin
					state<=1818;
					out<=161;
				end
				if(in == 4) begin
					state<=5707;
					out<=162;
				end
			end
			3719: begin
				if(in == 0) begin
					state<=3720;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=7609;
					out<=165;
				end
				if(in == 3) begin
					state<=1819;
					out<=166;
				end
				if(in == 4) begin
					state<=5708;
					out<=167;
				end
			end
			3720: begin
				if(in == 0) begin
					state<=3721;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=7610;
					out<=170;
				end
				if(in == 3) begin
					state<=1820;
					out<=171;
				end
				if(in == 4) begin
					state<=5709;
					out<=172;
				end
			end
			3721: begin
				if(in == 0) begin
					state<=3722;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=7611;
					out<=175;
				end
				if(in == 3) begin
					state<=1821;
					out<=176;
				end
				if(in == 4) begin
					state<=5710;
					out<=177;
				end
			end
			3722: begin
				if(in == 0) begin
					state<=3723;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=7612;
					out<=180;
				end
				if(in == 3) begin
					state<=1822;
					out<=181;
				end
				if(in == 4) begin
					state<=5711;
					out<=182;
				end
			end
			3723: begin
				if(in == 0) begin
					state<=3724;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=7613;
					out<=185;
				end
				if(in == 3) begin
					state<=1823;
					out<=186;
				end
				if(in == 4) begin
					state<=5712;
					out<=187;
				end
			end
			3724: begin
				if(in == 0) begin
					state<=3725;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=7614;
					out<=190;
				end
				if(in == 3) begin
					state<=1824;
					out<=191;
				end
				if(in == 4) begin
					state<=5713;
					out<=192;
				end
			end
			3725: begin
				if(in == 0) begin
					state<=3726;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=7615;
					out<=195;
				end
				if(in == 3) begin
					state<=1825;
					out<=196;
				end
				if(in == 4) begin
					state<=5714;
					out<=197;
				end
			end
			3726: begin
				if(in == 0) begin
					state<=3727;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=7616;
					out<=200;
				end
				if(in == 3) begin
					state<=1826;
					out<=201;
				end
				if(in == 4) begin
					state<=5715;
					out<=202;
				end
			end
			3727: begin
				if(in == 0) begin
					state<=3728;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=7617;
					out<=205;
				end
				if(in == 3) begin
					state<=1827;
					out<=206;
				end
				if(in == 4) begin
					state<=5716;
					out<=207;
				end
			end
			3728: begin
				if(in == 0) begin
					state<=3729;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=7618;
					out<=210;
				end
				if(in == 3) begin
					state<=1828;
					out<=211;
				end
				if(in == 4) begin
					state<=5717;
					out<=212;
				end
			end
			3729: begin
				if(in == 0) begin
					state<=3730;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=7619;
					out<=215;
				end
				if(in == 3) begin
					state<=1829;
					out<=216;
				end
				if(in == 4) begin
					state<=5718;
					out<=217;
				end
			end
			3730: begin
				if(in == 0) begin
					state<=3731;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=7620;
					out<=220;
				end
				if(in == 3) begin
					state<=1830;
					out<=221;
				end
				if(in == 4) begin
					state<=5719;
					out<=222;
				end
			end
			3731: begin
				if(in == 0) begin
					state<=3732;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=7621;
					out<=225;
				end
				if(in == 3) begin
					state<=1831;
					out<=226;
				end
				if(in == 4) begin
					state<=5720;
					out<=227;
				end
			end
			3732: begin
				if(in == 0) begin
					state<=3733;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=7622;
					out<=230;
				end
				if(in == 3) begin
					state<=1832;
					out<=231;
				end
				if(in == 4) begin
					state<=5721;
					out<=232;
				end
			end
			3733: begin
				if(in == 0) begin
					state<=3734;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=7623;
					out<=235;
				end
				if(in == 3) begin
					state<=1833;
					out<=236;
				end
				if(in == 4) begin
					state<=5722;
					out<=237;
				end
			end
			3734: begin
				if(in == 0) begin
					state<=3735;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=7624;
					out<=240;
				end
				if(in == 3) begin
					state<=1834;
					out<=241;
				end
				if(in == 4) begin
					state<=5723;
					out<=242;
				end
			end
			3735: begin
				if(in == 0) begin
					state<=3736;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=7625;
					out<=245;
				end
				if(in == 3) begin
					state<=1835;
					out<=246;
				end
				if(in == 4) begin
					state<=5724;
					out<=247;
				end
			end
			3736: begin
				if(in == 0) begin
					state<=3737;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=7626;
					out<=250;
				end
				if(in == 3) begin
					state<=1836;
					out<=251;
				end
				if(in == 4) begin
					state<=5725;
					out<=252;
				end
			end
			3737: begin
				if(in == 0) begin
					state<=3738;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=7627;
					out<=255;
				end
				if(in == 3) begin
					state<=1837;
					out<=0;
				end
				if(in == 4) begin
					state<=5726;
					out<=1;
				end
			end
			3738: begin
				if(in == 0) begin
					state<=3739;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=7628;
					out<=4;
				end
				if(in == 3) begin
					state<=1838;
					out<=5;
				end
				if(in == 4) begin
					state<=5727;
					out<=6;
				end
			end
			3739: begin
				if(in == 0) begin
					state<=3740;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=7629;
					out<=9;
				end
				if(in == 3) begin
					state<=1839;
					out<=10;
				end
				if(in == 4) begin
					state<=5728;
					out<=11;
				end
			end
			3740: begin
				if(in == 0) begin
					state<=3741;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=7630;
					out<=14;
				end
				if(in == 3) begin
					state<=1840;
					out<=15;
				end
				if(in == 4) begin
					state<=5729;
					out<=16;
				end
			end
			3741: begin
				if(in == 0) begin
					state<=3742;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=7631;
					out<=19;
				end
				if(in == 3) begin
					state<=1841;
					out<=20;
				end
				if(in == 4) begin
					state<=5730;
					out<=21;
				end
			end
			3742: begin
				if(in == 0) begin
					state<=3743;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=7632;
					out<=24;
				end
				if(in == 3) begin
					state<=1842;
					out<=25;
				end
				if(in == 4) begin
					state<=5731;
					out<=26;
				end
			end
			3743: begin
				if(in == 0) begin
					state<=3744;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=7633;
					out<=29;
				end
				if(in == 3) begin
					state<=1843;
					out<=30;
				end
				if(in == 4) begin
					state<=5732;
					out<=31;
				end
			end
			3744: begin
				if(in == 0) begin
					state<=3745;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=7634;
					out<=34;
				end
				if(in == 3) begin
					state<=1844;
					out<=35;
				end
				if(in == 4) begin
					state<=5733;
					out<=36;
				end
			end
			3745: begin
				if(in == 0) begin
					state<=3746;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=7635;
					out<=39;
				end
				if(in == 3) begin
					state<=1845;
					out<=40;
				end
				if(in == 4) begin
					state<=5734;
					out<=41;
				end
			end
			3746: begin
				if(in == 0) begin
					state<=3747;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=7636;
					out<=44;
				end
				if(in == 3) begin
					state<=1846;
					out<=45;
				end
				if(in == 4) begin
					state<=5735;
					out<=46;
				end
			end
			3747: begin
				if(in == 0) begin
					state<=3748;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=7637;
					out<=49;
				end
				if(in == 3) begin
					state<=1847;
					out<=50;
				end
				if(in == 4) begin
					state<=5736;
					out<=51;
				end
			end
			3748: begin
				if(in == 0) begin
					state<=3749;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=7638;
					out<=54;
				end
				if(in == 3) begin
					state<=1848;
					out<=55;
				end
				if(in == 4) begin
					state<=5737;
					out<=56;
				end
			end
			3749: begin
				if(in == 0) begin
					state<=3750;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=7639;
					out<=59;
				end
				if(in == 3) begin
					state<=1849;
					out<=60;
				end
				if(in == 4) begin
					state<=5738;
					out<=61;
				end
			end
			3750: begin
				if(in == 0) begin
					state<=3751;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=7640;
					out<=64;
				end
				if(in == 3) begin
					state<=1850;
					out<=65;
				end
				if(in == 4) begin
					state<=5739;
					out<=66;
				end
			end
			3751: begin
				if(in == 0) begin
					state<=3752;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=7641;
					out<=69;
				end
				if(in == 3) begin
					state<=1851;
					out<=70;
				end
				if(in == 4) begin
					state<=5740;
					out<=71;
				end
			end
			3752: begin
				if(in == 0) begin
					state<=3753;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=7642;
					out<=74;
				end
				if(in == 3) begin
					state<=1852;
					out<=75;
				end
				if(in == 4) begin
					state<=5741;
					out<=76;
				end
			end
			3753: begin
				if(in == 0) begin
					state<=3754;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=7643;
					out<=79;
				end
				if(in == 3) begin
					state<=1853;
					out<=80;
				end
				if(in == 4) begin
					state<=5742;
					out<=81;
				end
			end
			3754: begin
				if(in == 0) begin
					state<=3755;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=7644;
					out<=84;
				end
				if(in == 3) begin
					state<=1854;
					out<=85;
				end
				if(in == 4) begin
					state<=5743;
					out<=86;
				end
			end
			3755: begin
				if(in == 0) begin
					state<=3756;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=7645;
					out<=89;
				end
				if(in == 3) begin
					state<=1855;
					out<=90;
				end
				if(in == 4) begin
					state<=5744;
					out<=91;
				end
			end
			3756: begin
				if(in == 0) begin
					state<=3757;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=7646;
					out<=94;
				end
				if(in == 3) begin
					state<=1856;
					out<=95;
				end
				if(in == 4) begin
					state<=5745;
					out<=96;
				end
			end
			3757: begin
				if(in == 0) begin
					state<=3758;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=7647;
					out<=99;
				end
				if(in == 3) begin
					state<=1857;
					out<=100;
				end
				if(in == 4) begin
					state<=5746;
					out<=101;
				end
			end
			3758: begin
				if(in == 0) begin
					state<=3759;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=7648;
					out<=104;
				end
				if(in == 3) begin
					state<=1858;
					out<=105;
				end
				if(in == 4) begin
					state<=5747;
					out<=106;
				end
			end
			3759: begin
				if(in == 0) begin
					state<=3760;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=7649;
					out<=109;
				end
				if(in == 3) begin
					state<=1859;
					out<=110;
				end
				if(in == 4) begin
					state<=5748;
					out<=111;
				end
			end
			3760: begin
				if(in == 0) begin
					state<=3761;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=7650;
					out<=114;
				end
				if(in == 3) begin
					state<=1860;
					out<=115;
				end
				if(in == 4) begin
					state<=5749;
					out<=116;
				end
			end
			3761: begin
				if(in == 0) begin
					state<=3762;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=7651;
					out<=119;
				end
				if(in == 3) begin
					state<=1861;
					out<=120;
				end
				if(in == 4) begin
					state<=5750;
					out<=121;
				end
			end
			3762: begin
				if(in == 0) begin
					state<=3763;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=7652;
					out<=124;
				end
				if(in == 3) begin
					state<=1862;
					out<=125;
				end
				if(in == 4) begin
					state<=5751;
					out<=126;
				end
			end
			3763: begin
				if(in == 0) begin
					state<=3764;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=7653;
					out<=129;
				end
				if(in == 3) begin
					state<=1863;
					out<=130;
				end
				if(in == 4) begin
					state<=5752;
					out<=131;
				end
			end
			3764: begin
				if(in == 0) begin
					state<=3765;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=7654;
					out<=134;
				end
				if(in == 3) begin
					state<=1864;
					out<=135;
				end
				if(in == 4) begin
					state<=5753;
					out<=136;
				end
			end
			3765: begin
				if(in == 0) begin
					state<=3766;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=7655;
					out<=139;
				end
				if(in == 3) begin
					state<=1865;
					out<=140;
				end
				if(in == 4) begin
					state<=5754;
					out<=141;
				end
			end
			3766: begin
				if(in == 0) begin
					state<=3767;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=7656;
					out<=144;
				end
				if(in == 3) begin
					state<=1866;
					out<=145;
				end
				if(in == 4) begin
					state<=5755;
					out<=146;
				end
			end
			3767: begin
				if(in == 0) begin
					state<=3768;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=7657;
					out<=149;
				end
				if(in == 3) begin
					state<=1867;
					out<=150;
				end
				if(in == 4) begin
					state<=5756;
					out<=151;
				end
			end
			3768: begin
				if(in == 0) begin
					state<=3769;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=7658;
					out<=154;
				end
				if(in == 3) begin
					state<=1868;
					out<=155;
				end
				if(in == 4) begin
					state<=5757;
					out<=156;
				end
			end
			3769: begin
				if(in == 0) begin
					state<=3770;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=7659;
					out<=159;
				end
				if(in == 3) begin
					state<=1869;
					out<=160;
				end
				if(in == 4) begin
					state<=5758;
					out<=161;
				end
			end
			3770: begin
				if(in == 0) begin
					state<=3771;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=7660;
					out<=164;
				end
				if(in == 3) begin
					state<=1870;
					out<=165;
				end
				if(in == 4) begin
					state<=5759;
					out<=166;
				end
			end
			3771: begin
				if(in == 0) begin
					state<=3772;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=7661;
					out<=169;
				end
				if(in == 3) begin
					state<=1871;
					out<=170;
				end
				if(in == 4) begin
					state<=5760;
					out<=171;
				end
			end
			3772: begin
				if(in == 0) begin
					state<=3773;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=7662;
					out<=174;
				end
				if(in == 3) begin
					state<=1872;
					out<=175;
				end
				if(in == 4) begin
					state<=5761;
					out<=176;
				end
			end
			3773: begin
				if(in == 0) begin
					state<=3774;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=7663;
					out<=179;
				end
				if(in == 3) begin
					state<=1873;
					out<=180;
				end
				if(in == 4) begin
					state<=5762;
					out<=181;
				end
			end
			3774: begin
				if(in == 0) begin
					state<=3775;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=7664;
					out<=184;
				end
				if(in == 3) begin
					state<=1874;
					out<=185;
				end
				if(in == 4) begin
					state<=5763;
					out<=186;
				end
			end
			3775: begin
				if(in == 0) begin
					state<=3776;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=7665;
					out<=189;
				end
				if(in == 3) begin
					state<=1875;
					out<=190;
				end
				if(in == 4) begin
					state<=5764;
					out<=191;
				end
			end
			3776: begin
				if(in == 0) begin
					state<=3777;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=7666;
					out<=194;
				end
				if(in == 3) begin
					state<=1876;
					out<=195;
				end
				if(in == 4) begin
					state<=5765;
					out<=196;
				end
			end
			3777: begin
				if(in == 0) begin
					state<=3778;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=7667;
					out<=199;
				end
				if(in == 3) begin
					state<=1877;
					out<=200;
				end
				if(in == 4) begin
					state<=5766;
					out<=201;
				end
			end
			3778: begin
				if(in == 0) begin
					state<=3779;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=7668;
					out<=204;
				end
				if(in == 3) begin
					state<=1878;
					out<=205;
				end
				if(in == 4) begin
					state<=5767;
					out<=206;
				end
			end
			3779: begin
				if(in == 0) begin
					state<=3780;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=7669;
					out<=209;
				end
				if(in == 3) begin
					state<=1879;
					out<=210;
				end
				if(in == 4) begin
					state<=5768;
					out<=211;
				end
			end
			3780: begin
				if(in == 0) begin
					state<=3781;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=7670;
					out<=214;
				end
				if(in == 3) begin
					state<=1880;
					out<=215;
				end
				if(in == 4) begin
					state<=5769;
					out<=216;
				end
			end
			3781: begin
				if(in == 0) begin
					state<=3782;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=7671;
					out<=219;
				end
				if(in == 3) begin
					state<=1881;
					out<=220;
				end
				if(in == 4) begin
					state<=5770;
					out<=221;
				end
			end
			3782: begin
				if(in == 0) begin
					state<=3783;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=7672;
					out<=224;
				end
				if(in == 3) begin
					state<=1882;
					out<=225;
				end
				if(in == 4) begin
					state<=5771;
					out<=226;
				end
			end
			3783: begin
				if(in == 0) begin
					state<=3784;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=7673;
					out<=229;
				end
				if(in == 3) begin
					state<=1883;
					out<=230;
				end
				if(in == 4) begin
					state<=5772;
					out<=231;
				end
			end
			3784: begin
				if(in == 0) begin
					state<=3785;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=7674;
					out<=234;
				end
				if(in == 3) begin
					state<=1884;
					out<=235;
				end
				if(in == 4) begin
					state<=5773;
					out<=236;
				end
			end
			3785: begin
				if(in == 0) begin
					state<=3786;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=7675;
					out<=239;
				end
				if(in == 3) begin
					state<=1885;
					out<=240;
				end
				if(in == 4) begin
					state<=5774;
					out<=241;
				end
			end
			3786: begin
				if(in == 0) begin
					state<=3787;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=7676;
					out<=244;
				end
				if(in == 3) begin
					state<=1886;
					out<=245;
				end
				if(in == 4) begin
					state<=5775;
					out<=246;
				end
			end
			3787: begin
				if(in == 0) begin
					state<=3788;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=7677;
					out<=249;
				end
				if(in == 3) begin
					state<=1887;
					out<=250;
				end
				if(in == 4) begin
					state<=5776;
					out<=251;
				end
			end
			3788: begin
				if(in == 0) begin
					state<=3789;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=7678;
					out<=254;
				end
				if(in == 3) begin
					state<=1888;
					out<=255;
				end
				if(in == 4) begin
					state<=5777;
					out<=0;
				end
			end
			3789: begin
				if(in == 0) begin
					state<=3790;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=7679;
					out<=3;
				end
				if(in == 3) begin
					state<=1889;
					out<=4;
				end
				if(in == 4) begin
					state<=5778;
					out<=5;
				end
			end
			3790: begin
				if(in == 0) begin
					state<=3791;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=7680;
					out<=8;
				end
				if(in == 3) begin
					state<=1890;
					out<=9;
				end
				if(in == 4) begin
					state<=5779;
					out<=10;
				end
			end
			3791: begin
				if(in == 0) begin
					state<=3792;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=7681;
					out<=13;
				end
				if(in == 3) begin
					state<=1891;
					out<=14;
				end
				if(in == 4) begin
					state<=5780;
					out<=15;
				end
			end
			3792: begin
				if(in == 0) begin
					state<=3793;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=7682;
					out<=18;
				end
				if(in == 3) begin
					state<=1892;
					out<=19;
				end
				if(in == 4) begin
					state<=5781;
					out<=20;
				end
			end
			3793: begin
				if(in == 0) begin
					state<=3794;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=7683;
					out<=23;
				end
				if(in == 3) begin
					state<=1893;
					out<=24;
				end
				if(in == 4) begin
					state<=5782;
					out<=25;
				end
			end
			3794: begin
				if(in == 0) begin
					state<=3795;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=7684;
					out<=28;
				end
				if(in == 3) begin
					state<=1894;
					out<=29;
				end
				if(in == 4) begin
					state<=5783;
					out<=30;
				end
			end
			3795: begin
				if(in == 0) begin
					state<=3796;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=7685;
					out<=33;
				end
				if(in == 3) begin
					state<=1895;
					out<=34;
				end
				if(in == 4) begin
					state<=5784;
					out<=35;
				end
			end
			3796: begin
				if(in == 0) begin
					state<=3797;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=7686;
					out<=38;
				end
				if(in == 3) begin
					state<=1896;
					out<=39;
				end
				if(in == 4) begin
					state<=5785;
					out<=40;
				end
			end
			3797: begin
				if(in == 0) begin
					state<=3798;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=7687;
					out<=43;
				end
				if(in == 3) begin
					state<=1897;
					out<=44;
				end
				if(in == 4) begin
					state<=5786;
					out<=45;
				end
			end
			3798: begin
				if(in == 0) begin
					state<=3799;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=7688;
					out<=48;
				end
				if(in == 3) begin
					state<=1898;
					out<=49;
				end
				if(in == 4) begin
					state<=5787;
					out<=50;
				end
			end
			3799: begin
				if(in == 0) begin
					state<=3800;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=7689;
					out<=53;
				end
				if(in == 3) begin
					state<=1899;
					out<=54;
				end
				if(in == 4) begin
					state<=5788;
					out<=55;
				end
			end
			3800: begin
				if(in == 0) begin
					state<=3801;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=7690;
					out<=58;
				end
				if(in == 3) begin
					state<=1900;
					out<=59;
				end
				if(in == 4) begin
					state<=5789;
					out<=60;
				end
			end
			3801: begin
				if(in == 0) begin
					state<=3802;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=7691;
					out<=63;
				end
				if(in == 3) begin
					state<=1901;
					out<=64;
				end
				if(in == 4) begin
					state<=5790;
					out<=65;
				end
			end
			3802: begin
				if(in == 0) begin
					state<=3803;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=7692;
					out<=68;
				end
				if(in == 3) begin
					state<=1902;
					out<=69;
				end
				if(in == 4) begin
					state<=5791;
					out<=70;
				end
			end
			3803: begin
				if(in == 0) begin
					state<=3804;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=7693;
					out<=73;
				end
				if(in == 3) begin
					state<=1903;
					out<=74;
				end
				if(in == 4) begin
					state<=5792;
					out<=75;
				end
			end
			3804: begin
				if(in == 0) begin
					state<=3805;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=7694;
					out<=78;
				end
				if(in == 3) begin
					state<=1904;
					out<=79;
				end
				if(in == 4) begin
					state<=5793;
					out<=80;
				end
			end
			3805: begin
				if(in == 0) begin
					state<=3806;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=7695;
					out<=83;
				end
				if(in == 3) begin
					state<=1905;
					out<=84;
				end
				if(in == 4) begin
					state<=5794;
					out<=85;
				end
			end
			3806: begin
				if(in == 0) begin
					state<=3807;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=7696;
					out<=88;
				end
				if(in == 3) begin
					state<=1906;
					out<=89;
				end
				if(in == 4) begin
					state<=5795;
					out<=90;
				end
			end
			3807: begin
				if(in == 0) begin
					state<=3808;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=7697;
					out<=93;
				end
				if(in == 3) begin
					state<=1907;
					out<=94;
				end
				if(in == 4) begin
					state<=5796;
					out<=95;
				end
			end
			3808: begin
				if(in == 0) begin
					state<=3809;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=7698;
					out<=98;
				end
				if(in == 3) begin
					state<=1908;
					out<=99;
				end
				if(in == 4) begin
					state<=5797;
					out<=100;
				end
			end
			3809: begin
				if(in == 0) begin
					state<=3810;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=7699;
					out<=103;
				end
				if(in == 3) begin
					state<=1909;
					out<=104;
				end
				if(in == 4) begin
					state<=5798;
					out<=105;
				end
			end
			3810: begin
				if(in == 0) begin
					state<=3811;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=7700;
					out<=108;
				end
				if(in == 3) begin
					state<=1910;
					out<=109;
				end
				if(in == 4) begin
					state<=5799;
					out<=110;
				end
			end
			3811: begin
				if(in == 0) begin
					state<=3812;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=7701;
					out<=113;
				end
				if(in == 3) begin
					state<=1911;
					out<=114;
				end
				if(in == 4) begin
					state<=5800;
					out<=115;
				end
			end
			3812: begin
				if(in == 0) begin
					state<=3813;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=7702;
					out<=118;
				end
				if(in == 3) begin
					state<=1912;
					out<=119;
				end
				if(in == 4) begin
					state<=5801;
					out<=120;
				end
			end
			3813: begin
				if(in == 0) begin
					state<=3814;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=7703;
					out<=123;
				end
				if(in == 3) begin
					state<=1913;
					out<=124;
				end
				if(in == 4) begin
					state<=5802;
					out<=125;
				end
			end
			3814: begin
				if(in == 0) begin
					state<=3815;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=7704;
					out<=128;
				end
				if(in == 3) begin
					state<=1914;
					out<=129;
				end
				if(in == 4) begin
					state<=5803;
					out<=130;
				end
			end
			3815: begin
				if(in == 0) begin
					state<=3816;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=7705;
					out<=133;
				end
				if(in == 3) begin
					state<=1915;
					out<=134;
				end
				if(in == 4) begin
					state<=5804;
					out<=135;
				end
			end
			3816: begin
				if(in == 0) begin
					state<=3817;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=7706;
					out<=138;
				end
				if(in == 3) begin
					state<=1916;
					out<=139;
				end
				if(in == 4) begin
					state<=5805;
					out<=140;
				end
			end
			3817: begin
				if(in == 0) begin
					state<=3818;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=7707;
					out<=143;
				end
				if(in == 3) begin
					state<=1917;
					out<=144;
				end
				if(in == 4) begin
					state<=5806;
					out<=145;
				end
			end
			3818: begin
				if(in == 0) begin
					state<=3819;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=7708;
					out<=148;
				end
				if(in == 3) begin
					state<=1918;
					out<=149;
				end
				if(in == 4) begin
					state<=5807;
					out<=150;
				end
			end
			3819: begin
				if(in == 0) begin
					state<=3820;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=7709;
					out<=153;
				end
				if(in == 3) begin
					state<=1919;
					out<=154;
				end
				if(in == 4) begin
					state<=5808;
					out<=155;
				end
			end
			3820: begin
				if(in == 0) begin
					state<=3821;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=7710;
					out<=158;
				end
				if(in == 3) begin
					state<=1920;
					out<=159;
				end
				if(in == 4) begin
					state<=5809;
					out<=160;
				end
			end
			3821: begin
				if(in == 0) begin
					state<=3822;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=7711;
					out<=163;
				end
				if(in == 3) begin
					state<=1921;
					out<=164;
				end
				if(in == 4) begin
					state<=5810;
					out<=165;
				end
			end
			3822: begin
				if(in == 0) begin
					state<=3823;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=7712;
					out<=168;
				end
				if(in == 3) begin
					state<=1922;
					out<=169;
				end
				if(in == 4) begin
					state<=5811;
					out<=170;
				end
			end
			3823: begin
				if(in == 0) begin
					state<=3824;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=7713;
					out<=173;
				end
				if(in == 3) begin
					state<=1923;
					out<=174;
				end
				if(in == 4) begin
					state<=5812;
					out<=175;
				end
			end
			3824: begin
				if(in == 0) begin
					state<=3825;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=7714;
					out<=178;
				end
				if(in == 3) begin
					state<=1924;
					out<=179;
				end
				if(in == 4) begin
					state<=5813;
					out<=180;
				end
			end
			3825: begin
				if(in == 0) begin
					state<=3826;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=7715;
					out<=183;
				end
				if(in == 3) begin
					state<=1925;
					out<=184;
				end
				if(in == 4) begin
					state<=5814;
					out<=185;
				end
			end
			3826: begin
				if(in == 0) begin
					state<=3827;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=7716;
					out<=188;
				end
				if(in == 3) begin
					state<=1926;
					out<=189;
				end
				if(in == 4) begin
					state<=5815;
					out<=190;
				end
			end
			3827: begin
				if(in == 0) begin
					state<=3828;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=7717;
					out<=193;
				end
				if(in == 3) begin
					state<=1927;
					out<=194;
				end
				if(in == 4) begin
					state<=5816;
					out<=195;
				end
			end
			3828: begin
				if(in == 0) begin
					state<=3829;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=7718;
					out<=198;
				end
				if(in == 3) begin
					state<=1928;
					out<=199;
				end
				if(in == 4) begin
					state<=5817;
					out<=200;
				end
			end
			3829: begin
				if(in == 0) begin
					state<=3830;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=7719;
					out<=203;
				end
				if(in == 3) begin
					state<=1929;
					out<=204;
				end
				if(in == 4) begin
					state<=5818;
					out<=205;
				end
			end
			3830: begin
				if(in == 0) begin
					state<=3831;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=7720;
					out<=208;
				end
				if(in == 3) begin
					state<=1930;
					out<=209;
				end
				if(in == 4) begin
					state<=5819;
					out<=210;
				end
			end
			3831: begin
				if(in == 0) begin
					state<=3832;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=7721;
					out<=213;
				end
				if(in == 3) begin
					state<=1931;
					out<=214;
				end
				if(in == 4) begin
					state<=5820;
					out<=215;
				end
			end
			3832: begin
				if(in == 0) begin
					state<=3833;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=7722;
					out<=218;
				end
				if(in == 3) begin
					state<=1932;
					out<=219;
				end
				if(in == 4) begin
					state<=5821;
					out<=220;
				end
			end
			3833: begin
				if(in == 0) begin
					state<=3834;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=7723;
					out<=223;
				end
				if(in == 3) begin
					state<=1933;
					out<=224;
				end
				if(in == 4) begin
					state<=5822;
					out<=225;
				end
			end
			3834: begin
				if(in == 0) begin
					state<=3835;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=7724;
					out<=228;
				end
				if(in == 3) begin
					state<=1934;
					out<=229;
				end
				if(in == 4) begin
					state<=5823;
					out<=230;
				end
			end
			3835: begin
				if(in == 0) begin
					state<=3836;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=7725;
					out<=233;
				end
				if(in == 3) begin
					state<=1935;
					out<=234;
				end
				if(in == 4) begin
					state<=5824;
					out<=235;
				end
			end
			3836: begin
				if(in == 0) begin
					state<=3837;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=7726;
					out<=238;
				end
				if(in == 3) begin
					state<=1936;
					out<=239;
				end
				if(in == 4) begin
					state<=5825;
					out<=240;
				end
			end
			3837: begin
				if(in == 0) begin
					state<=3838;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=7727;
					out<=243;
				end
				if(in == 3) begin
					state<=1937;
					out<=244;
				end
				if(in == 4) begin
					state<=5826;
					out<=245;
				end
			end
			3838: begin
				if(in == 0) begin
					state<=3839;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=7728;
					out<=248;
				end
				if(in == 3) begin
					state<=1938;
					out<=249;
				end
				if(in == 4) begin
					state<=5827;
					out<=250;
				end
			end
			3839: begin
				if(in == 0) begin
					state<=3840;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=7729;
					out<=253;
				end
				if(in == 3) begin
					state<=1939;
					out<=254;
				end
				if(in == 4) begin
					state<=5828;
					out<=255;
				end
			end
			3840: begin
				if(in == 0) begin
					state<=3841;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=7730;
					out<=2;
				end
				if(in == 3) begin
					state<=1940;
					out<=3;
				end
				if(in == 4) begin
					state<=5829;
					out<=4;
				end
			end
			3841: begin
				if(in == 0) begin
					state<=3842;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=7731;
					out<=7;
				end
				if(in == 3) begin
					state<=1941;
					out<=8;
				end
				if(in == 4) begin
					state<=5830;
					out<=9;
				end
			end
			3842: begin
				if(in == 0) begin
					state<=3843;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=7732;
					out<=12;
				end
				if(in == 3) begin
					state<=1942;
					out<=13;
				end
				if(in == 4) begin
					state<=5831;
					out<=14;
				end
			end
			3843: begin
				if(in == 0) begin
					state<=3844;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=7733;
					out<=17;
				end
				if(in == 3) begin
					state<=1943;
					out<=18;
				end
				if(in == 4) begin
					state<=5832;
					out<=19;
				end
			end
			3844: begin
				if(in == 0) begin
					state<=3845;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=7734;
					out<=22;
				end
				if(in == 3) begin
					state<=1944;
					out<=23;
				end
				if(in == 4) begin
					state<=5833;
					out<=24;
				end
			end
			3845: begin
				if(in == 0) begin
					state<=3846;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=7735;
					out<=27;
				end
				if(in == 3) begin
					state<=1945;
					out<=28;
				end
				if(in == 4) begin
					state<=5834;
					out<=29;
				end
			end
			3846: begin
				if(in == 0) begin
					state<=3847;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=7736;
					out<=32;
				end
				if(in == 3) begin
					state<=1946;
					out<=33;
				end
				if(in == 4) begin
					state<=5835;
					out<=34;
				end
			end
			3847: begin
				if(in == 0) begin
					state<=3848;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=7737;
					out<=37;
				end
				if(in == 3) begin
					state<=1947;
					out<=38;
				end
				if(in == 4) begin
					state<=5836;
					out<=39;
				end
			end
			3848: begin
				if(in == 0) begin
					state<=3849;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=7738;
					out<=42;
				end
				if(in == 3) begin
					state<=1948;
					out<=43;
				end
				if(in == 4) begin
					state<=5837;
					out<=44;
				end
			end
			3849: begin
				if(in == 0) begin
					state<=3850;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=7739;
					out<=47;
				end
				if(in == 3) begin
					state<=1949;
					out<=48;
				end
				if(in == 4) begin
					state<=5838;
					out<=49;
				end
			end
			3850: begin
				if(in == 0) begin
					state<=3851;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=7740;
					out<=52;
				end
				if(in == 3) begin
					state<=1950;
					out<=53;
				end
				if(in == 4) begin
					state<=5839;
					out<=54;
				end
			end
			3851: begin
				if(in == 0) begin
					state<=3852;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=7741;
					out<=57;
				end
				if(in == 3) begin
					state<=1951;
					out<=58;
				end
				if(in == 4) begin
					state<=5840;
					out<=59;
				end
			end
			3852: begin
				if(in == 0) begin
					state<=3853;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=7742;
					out<=62;
				end
				if(in == 3) begin
					state<=1952;
					out<=63;
				end
				if(in == 4) begin
					state<=5841;
					out<=64;
				end
			end
			3853: begin
				if(in == 0) begin
					state<=3854;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=7743;
					out<=67;
				end
				if(in == 3) begin
					state<=1953;
					out<=68;
				end
				if(in == 4) begin
					state<=5842;
					out<=69;
				end
			end
			3854: begin
				if(in == 0) begin
					state<=3855;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=7744;
					out<=72;
				end
				if(in == 3) begin
					state<=1954;
					out<=73;
				end
				if(in == 4) begin
					state<=5843;
					out<=74;
				end
			end
			3855: begin
				if(in == 0) begin
					state<=3856;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=7745;
					out<=77;
				end
				if(in == 3) begin
					state<=1955;
					out<=78;
				end
				if(in == 4) begin
					state<=5844;
					out<=79;
				end
			end
			3856: begin
				if(in == 0) begin
					state<=3857;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=7746;
					out<=82;
				end
				if(in == 3) begin
					state<=1956;
					out<=83;
				end
				if(in == 4) begin
					state<=5845;
					out<=84;
				end
			end
			3857: begin
				if(in == 0) begin
					state<=3858;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=7747;
					out<=87;
				end
				if(in == 3) begin
					state<=1957;
					out<=88;
				end
				if(in == 4) begin
					state<=5846;
					out<=89;
				end
			end
			3858: begin
				if(in == 0) begin
					state<=3859;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=7748;
					out<=92;
				end
				if(in == 3) begin
					state<=1958;
					out<=93;
				end
				if(in == 4) begin
					state<=5847;
					out<=94;
				end
			end
			3859: begin
				if(in == 0) begin
					state<=3860;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=7749;
					out<=97;
				end
				if(in == 3) begin
					state<=1959;
					out<=98;
				end
				if(in == 4) begin
					state<=5848;
					out<=99;
				end
			end
			3860: begin
				if(in == 0) begin
					state<=3861;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=7750;
					out<=102;
				end
				if(in == 3) begin
					state<=1960;
					out<=103;
				end
				if(in == 4) begin
					state<=5849;
					out<=104;
				end
			end
			3861: begin
				if(in == 0) begin
					state<=3862;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=7751;
					out<=107;
				end
				if(in == 3) begin
					state<=1961;
					out<=108;
				end
				if(in == 4) begin
					state<=5850;
					out<=109;
				end
			end
			3862: begin
				if(in == 0) begin
					state<=3863;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=7752;
					out<=112;
				end
				if(in == 3) begin
					state<=1962;
					out<=113;
				end
				if(in == 4) begin
					state<=5851;
					out<=114;
				end
			end
			3863: begin
				if(in == 0) begin
					state<=3864;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=7753;
					out<=117;
				end
				if(in == 3) begin
					state<=1963;
					out<=118;
				end
				if(in == 4) begin
					state<=5852;
					out<=119;
				end
			end
			3864: begin
				if(in == 0) begin
					state<=3865;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=7754;
					out<=122;
				end
				if(in == 3) begin
					state<=1964;
					out<=123;
				end
				if(in == 4) begin
					state<=5853;
					out<=124;
				end
			end
			3865: begin
				if(in == 0) begin
					state<=3866;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=7755;
					out<=127;
				end
				if(in == 3) begin
					state<=1965;
					out<=128;
				end
				if(in == 4) begin
					state<=5854;
					out<=129;
				end
			end
			3866: begin
				if(in == 0) begin
					state<=3867;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=7756;
					out<=132;
				end
				if(in == 3) begin
					state<=1966;
					out<=133;
				end
				if(in == 4) begin
					state<=5855;
					out<=134;
				end
			end
			3867: begin
				if(in == 0) begin
					state<=3868;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=7757;
					out<=137;
				end
				if(in == 3) begin
					state<=1967;
					out<=138;
				end
				if(in == 4) begin
					state<=5856;
					out<=139;
				end
			end
			3868: begin
				if(in == 0) begin
					state<=3869;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=7758;
					out<=142;
				end
				if(in == 3) begin
					state<=1968;
					out<=143;
				end
				if(in == 4) begin
					state<=5857;
					out<=144;
				end
			end
			3869: begin
				if(in == 0) begin
					state<=3870;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=7759;
					out<=147;
				end
				if(in == 3) begin
					state<=1969;
					out<=148;
				end
				if(in == 4) begin
					state<=5858;
					out<=149;
				end
			end
			3870: begin
				if(in == 0) begin
					state<=3871;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=7760;
					out<=152;
				end
				if(in == 3) begin
					state<=1970;
					out<=153;
				end
				if(in == 4) begin
					state<=5859;
					out<=154;
				end
			end
			3871: begin
				if(in == 0) begin
					state<=3872;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=7761;
					out<=157;
				end
				if(in == 3) begin
					state<=1971;
					out<=158;
				end
				if(in == 4) begin
					state<=5860;
					out<=159;
				end
			end
			3872: begin
				if(in == 0) begin
					state<=3873;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=7762;
					out<=162;
				end
				if(in == 3) begin
					state<=1972;
					out<=163;
				end
				if(in == 4) begin
					state<=5861;
					out<=164;
				end
			end
			3873: begin
				if(in == 0) begin
					state<=3874;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=7763;
					out<=167;
				end
				if(in == 3) begin
					state<=1973;
					out<=168;
				end
				if(in == 4) begin
					state<=5862;
					out<=169;
				end
			end
			3874: begin
				if(in == 0) begin
					state<=3875;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=7764;
					out<=172;
				end
				if(in == 3) begin
					state<=1974;
					out<=173;
				end
				if(in == 4) begin
					state<=5863;
					out<=174;
				end
			end
			3875: begin
				if(in == 0) begin
					state<=3876;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=7765;
					out<=177;
				end
				if(in == 3) begin
					state<=1975;
					out<=178;
				end
				if(in == 4) begin
					state<=5864;
					out<=179;
				end
			end
			3876: begin
				if(in == 0) begin
					state<=3877;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=7766;
					out<=182;
				end
				if(in == 3) begin
					state<=1976;
					out<=183;
				end
				if(in == 4) begin
					state<=5865;
					out<=184;
				end
			end
			3877: begin
				if(in == 0) begin
					state<=3878;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=7767;
					out<=187;
				end
				if(in == 3) begin
					state<=1977;
					out<=188;
				end
				if(in == 4) begin
					state<=5866;
					out<=189;
				end
			end
			3878: begin
				if(in == 0) begin
					state<=3879;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=7768;
					out<=192;
				end
				if(in == 3) begin
					state<=1978;
					out<=193;
				end
				if(in == 4) begin
					state<=5867;
					out<=194;
				end
			end
			3879: begin
				if(in == 0) begin
					state<=3880;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=7769;
					out<=197;
				end
				if(in == 3) begin
					state<=1979;
					out<=198;
				end
				if(in == 4) begin
					state<=5868;
					out<=199;
				end
			end
			3880: begin
				if(in == 0) begin
					state<=3881;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=7770;
					out<=202;
				end
				if(in == 3) begin
					state<=1980;
					out<=203;
				end
				if(in == 4) begin
					state<=5869;
					out<=204;
				end
			end
			3881: begin
				if(in == 0) begin
					state<=3882;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=7771;
					out<=207;
				end
				if(in == 3) begin
					state<=1981;
					out<=208;
				end
				if(in == 4) begin
					state<=5870;
					out<=209;
				end
			end
			3882: begin
				if(in == 0) begin
					state<=3883;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=7772;
					out<=212;
				end
				if(in == 3) begin
					state<=1982;
					out<=213;
				end
				if(in == 4) begin
					state<=5871;
					out<=214;
				end
			end
			3883: begin
				if(in == 0) begin
					state<=3884;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=7773;
					out<=217;
				end
				if(in == 3) begin
					state<=1983;
					out<=218;
				end
				if(in == 4) begin
					state<=5872;
					out<=219;
				end
			end
			3884: begin
				if(in == 0) begin
					state<=3885;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=7774;
					out<=222;
				end
				if(in == 3) begin
					state<=1984;
					out<=223;
				end
				if(in == 4) begin
					state<=5873;
					out<=224;
				end
			end
			3885: begin
				if(in == 0) begin
					state<=3886;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=7775;
					out<=227;
				end
				if(in == 3) begin
					state<=1985;
					out<=228;
				end
				if(in == 4) begin
					state<=5874;
					out<=229;
				end
			end
			3886: begin
				if(in == 0) begin
					state<=3887;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=7776;
					out<=232;
				end
				if(in == 3) begin
					state<=1986;
					out<=233;
				end
				if(in == 4) begin
					state<=5875;
					out<=234;
				end
			end
			3887: begin
				if(in == 0) begin
					state<=3888;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=7777;
					out<=237;
				end
				if(in == 3) begin
					state<=1987;
					out<=238;
				end
				if(in == 4) begin
					state<=5876;
					out<=239;
				end
			end
			3888: begin
				if(in == 0) begin
					state<=3889;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=7778;
					out<=242;
				end
				if(in == 3) begin
					state<=1988;
					out<=243;
				end
				if(in == 4) begin
					state<=5877;
					out<=244;
				end
			end
			3889: begin
				if(in == 0) begin
					state<=3890;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=7779;
					out<=247;
				end
				if(in == 3) begin
					state<=1989;
					out<=248;
				end
				if(in == 4) begin
					state<=5878;
					out<=249;
				end
			end
			3890: begin
				if(in == 0) begin
					state<=3891;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=7780;
					out<=252;
				end
				if(in == 3) begin
					state<=1990;
					out<=253;
				end
				if(in == 4) begin
					state<=5879;
					out<=254;
				end
			end
			3891: begin
				if(in == 0) begin
					state<=3892;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=7781;
					out<=1;
				end
				if(in == 3) begin
					state<=1991;
					out<=2;
				end
				if(in == 4) begin
					state<=5880;
					out<=3;
				end
			end
			3892: begin
				if(in == 0) begin
					state<=3893;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=7782;
					out<=6;
				end
				if(in == 3) begin
					state<=1992;
					out<=7;
				end
				if(in == 4) begin
					state<=5881;
					out<=8;
				end
			end
			3893: begin
				if(in == 0) begin
					state<=3894;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=7783;
					out<=11;
				end
				if(in == 3) begin
					state<=1993;
					out<=12;
				end
				if(in == 4) begin
					state<=5882;
					out<=13;
				end
			end
			3894: begin
				if(in == 0) begin
					state<=3895;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=7784;
					out<=16;
				end
				if(in == 3) begin
					state<=1994;
					out<=17;
				end
				if(in == 4) begin
					state<=5883;
					out<=18;
				end
			end
			3895: begin
				if(in == 0) begin
					state<=3896;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=7785;
					out<=21;
				end
				if(in == 3) begin
					state<=1995;
					out<=22;
				end
				if(in == 4) begin
					state<=5884;
					out<=23;
				end
			end
			3896: begin
				if(in == 0) begin
					state<=3897;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=7786;
					out<=26;
				end
				if(in == 3) begin
					state<=1996;
					out<=27;
				end
				if(in == 4) begin
					state<=5885;
					out<=28;
				end
			end
			3897: begin
				if(in == 0) begin
					state<=3898;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=7787;
					out<=31;
				end
				if(in == 3) begin
					state<=1997;
					out<=32;
				end
				if(in == 4) begin
					state<=5886;
					out<=33;
				end
			end
			3898: begin
				if(in == 0) begin
					state<=2275;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=6164;
					out<=36;
				end
				if(in == 3) begin
					state<=1998;
					out<=37;
				end
				if(in == 4) begin
					state<=5887;
					out<=38;
				end
			end
			3899: begin
				if(in == 0) begin
					state<=3910;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=12;
					out<=41;
				end
				if(in == 3) begin
					state<=5899;
					out<=42;
				end
				if(in == 4) begin
					state<=2010;
					out<=43;
				end
			end
			3900: begin
				if(in == 0) begin
					state<=3911;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=13;
					out<=46;
				end
				if(in == 3) begin
					state<=5900;
					out<=47;
				end
				if(in == 4) begin
					state<=2011;
					out<=48;
				end
			end
			3901: begin
				if(in == 0) begin
					state<=3912;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=14;
					out<=51;
				end
				if(in == 3) begin
					state<=5901;
					out<=52;
				end
				if(in == 4) begin
					state<=2012;
					out<=53;
				end
			end
			3902: begin
				if(in == 0) begin
					state<=3913;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=15;
					out<=56;
				end
				if(in == 3) begin
					state<=5902;
					out<=57;
				end
				if(in == 4) begin
					state<=2013;
					out<=58;
				end
			end
			3903: begin
				if(in == 0) begin
					state<=3914;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=16;
					out<=61;
				end
				if(in == 3) begin
					state<=5903;
					out<=62;
				end
				if(in == 4) begin
					state<=2014;
					out<=63;
				end
			end
			3904: begin
				if(in == 0) begin
					state<=3915;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=17;
					out<=66;
				end
				if(in == 3) begin
					state<=5904;
					out<=67;
				end
				if(in == 4) begin
					state<=2015;
					out<=68;
				end
			end
			3905: begin
				if(in == 0) begin
					state<=3916;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=18;
					out<=71;
				end
				if(in == 3) begin
					state<=5905;
					out<=72;
				end
				if(in == 4) begin
					state<=2016;
					out<=73;
				end
			end
			3906: begin
				if(in == 0) begin
					state<=3917;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=19;
					out<=76;
				end
				if(in == 3) begin
					state<=5906;
					out<=77;
				end
				if(in == 4) begin
					state<=2017;
					out<=78;
				end
			end
			3907: begin
				if(in == 0) begin
					state<=3918;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=20;
					out<=81;
				end
				if(in == 3) begin
					state<=5907;
					out<=82;
				end
				if(in == 4) begin
					state<=2018;
					out<=83;
				end
			end
			3908: begin
				if(in == 0) begin
					state<=3909;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=11;
					out<=86;
				end
				if(in == 3) begin
					state<=5898;
					out<=87;
				end
				if(in == 4) begin
					state<=2009;
					out<=88;
				end
			end
			3909: begin
				if(in == 0) begin
					state<=3920;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=22;
					out<=91;
				end
				if(in == 3) begin
					state<=5909;
					out<=92;
				end
				if(in == 4) begin
					state<=2020;
					out<=93;
				end
			end
			3910: begin
				if(in == 0) begin
					state<=3921;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=23;
					out<=96;
				end
				if(in == 3) begin
					state<=5910;
					out<=97;
				end
				if(in == 4) begin
					state<=2021;
					out<=98;
				end
			end
			3911: begin
				if(in == 0) begin
					state<=3922;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=24;
					out<=101;
				end
				if(in == 3) begin
					state<=5911;
					out<=102;
				end
				if(in == 4) begin
					state<=2022;
					out<=103;
				end
			end
			3912: begin
				if(in == 0) begin
					state<=3923;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=25;
					out<=106;
				end
				if(in == 3) begin
					state<=5912;
					out<=107;
				end
				if(in == 4) begin
					state<=2023;
					out<=108;
				end
			end
			3913: begin
				if(in == 0) begin
					state<=3924;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=26;
					out<=111;
				end
				if(in == 3) begin
					state<=5913;
					out<=112;
				end
				if(in == 4) begin
					state<=2024;
					out<=113;
				end
			end
			3914: begin
				if(in == 0) begin
					state<=3925;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=27;
					out<=116;
				end
				if(in == 3) begin
					state<=5914;
					out<=117;
				end
				if(in == 4) begin
					state<=2025;
					out<=118;
				end
			end
			3915: begin
				if(in == 0) begin
					state<=3926;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=28;
					out<=121;
				end
				if(in == 3) begin
					state<=5915;
					out<=122;
				end
				if(in == 4) begin
					state<=2026;
					out<=123;
				end
			end
			3916: begin
				if(in == 0) begin
					state<=3927;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=29;
					out<=126;
				end
				if(in == 3) begin
					state<=5916;
					out<=127;
				end
				if(in == 4) begin
					state<=2027;
					out<=128;
				end
			end
			3917: begin
				if(in == 0) begin
					state<=3928;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=30;
					out<=131;
				end
				if(in == 3) begin
					state<=5917;
					out<=132;
				end
				if(in == 4) begin
					state<=2028;
					out<=133;
				end
			end
			3918: begin
				if(in == 0) begin
					state<=3919;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=21;
					out<=136;
				end
				if(in == 3) begin
					state<=5908;
					out<=137;
				end
				if(in == 4) begin
					state<=2019;
					out<=138;
				end
			end
			3919: begin
				if(in == 0) begin
					state<=3930;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=32;
					out<=141;
				end
				if(in == 3) begin
					state<=5919;
					out<=142;
				end
				if(in == 4) begin
					state<=2030;
					out<=143;
				end
			end
			3920: begin
				if(in == 0) begin
					state<=3931;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=33;
					out<=146;
				end
				if(in == 3) begin
					state<=5920;
					out<=147;
				end
				if(in == 4) begin
					state<=2031;
					out<=148;
				end
			end
			3921: begin
				if(in == 0) begin
					state<=3932;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=34;
					out<=151;
				end
				if(in == 3) begin
					state<=5921;
					out<=152;
				end
				if(in == 4) begin
					state<=2032;
					out<=153;
				end
			end
			3922: begin
				if(in == 0) begin
					state<=3933;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=35;
					out<=156;
				end
				if(in == 3) begin
					state<=5922;
					out<=157;
				end
				if(in == 4) begin
					state<=2033;
					out<=158;
				end
			end
			3923: begin
				if(in == 0) begin
					state<=3934;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=36;
					out<=161;
				end
				if(in == 3) begin
					state<=5923;
					out<=162;
				end
				if(in == 4) begin
					state<=2034;
					out<=163;
				end
			end
			3924: begin
				if(in == 0) begin
					state<=3935;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=37;
					out<=166;
				end
				if(in == 3) begin
					state<=5924;
					out<=167;
				end
				if(in == 4) begin
					state<=2035;
					out<=168;
				end
			end
			3925: begin
				if(in == 0) begin
					state<=3936;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=38;
					out<=171;
				end
				if(in == 3) begin
					state<=5925;
					out<=172;
				end
				if(in == 4) begin
					state<=2036;
					out<=173;
				end
			end
			3926: begin
				if(in == 0) begin
					state<=3937;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=39;
					out<=176;
				end
				if(in == 3) begin
					state<=5926;
					out<=177;
				end
				if(in == 4) begin
					state<=2037;
					out<=178;
				end
			end
			3927: begin
				if(in == 0) begin
					state<=3938;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=40;
					out<=181;
				end
				if(in == 3) begin
					state<=5927;
					out<=182;
				end
				if(in == 4) begin
					state<=2038;
					out<=183;
				end
			end
			3928: begin
				if(in == 0) begin
					state<=3929;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=31;
					out<=186;
				end
				if(in == 3) begin
					state<=5918;
					out<=187;
				end
				if(in == 4) begin
					state<=2029;
					out<=188;
				end
			end
			3929: begin
				if(in == 0) begin
					state<=3940;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=42;
					out<=191;
				end
				if(in == 3) begin
					state<=5929;
					out<=192;
				end
				if(in == 4) begin
					state<=2040;
					out<=193;
				end
			end
			3930: begin
				if(in == 0) begin
					state<=3941;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=43;
					out<=196;
				end
				if(in == 3) begin
					state<=5930;
					out<=197;
				end
				if(in == 4) begin
					state<=2041;
					out<=198;
				end
			end
			3931: begin
				if(in == 0) begin
					state<=3942;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=44;
					out<=201;
				end
				if(in == 3) begin
					state<=5931;
					out<=202;
				end
				if(in == 4) begin
					state<=2042;
					out<=203;
				end
			end
			3932: begin
				if(in == 0) begin
					state<=3943;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=45;
					out<=206;
				end
				if(in == 3) begin
					state<=5932;
					out<=207;
				end
				if(in == 4) begin
					state<=2043;
					out<=208;
				end
			end
			3933: begin
				if(in == 0) begin
					state<=3944;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=46;
					out<=211;
				end
				if(in == 3) begin
					state<=5933;
					out<=212;
				end
				if(in == 4) begin
					state<=2044;
					out<=213;
				end
			end
			3934: begin
				if(in == 0) begin
					state<=3945;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=47;
					out<=216;
				end
				if(in == 3) begin
					state<=5934;
					out<=217;
				end
				if(in == 4) begin
					state<=2045;
					out<=218;
				end
			end
			3935: begin
				if(in == 0) begin
					state<=3946;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=48;
					out<=221;
				end
				if(in == 3) begin
					state<=5935;
					out<=222;
				end
				if(in == 4) begin
					state<=2046;
					out<=223;
				end
			end
			3936: begin
				if(in == 0) begin
					state<=3947;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=49;
					out<=226;
				end
				if(in == 3) begin
					state<=5936;
					out<=227;
				end
				if(in == 4) begin
					state<=2047;
					out<=228;
				end
			end
			3937: begin
				if(in == 0) begin
					state<=3948;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=50;
					out<=231;
				end
				if(in == 3) begin
					state<=5937;
					out<=232;
				end
				if(in == 4) begin
					state<=2048;
					out<=233;
				end
			end
			3938: begin
				if(in == 0) begin
					state<=3939;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=41;
					out<=236;
				end
				if(in == 3) begin
					state<=5928;
					out<=237;
				end
				if(in == 4) begin
					state<=2039;
					out<=238;
				end
			end
			3939: begin
				if(in == 0) begin
					state<=5219;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=1330;
					out<=241;
				end
				if(in == 3) begin
					state<=7151;
					out<=242;
				end
				if(in == 4) begin
					state<=3262;
					out<=243;
				end
			end
			3940: begin
				if(in == 0) begin
					state<=5220;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=1331;
					out<=246;
				end
				if(in == 3) begin
					state<=7152;
					out<=247;
				end
				if(in == 4) begin
					state<=3263;
					out<=248;
				end
			end
			3941: begin
				if(in == 0) begin
					state<=5221;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=1332;
					out<=251;
				end
				if(in == 3) begin
					state<=7153;
					out<=252;
				end
				if(in == 4) begin
					state<=3264;
					out<=253;
				end
			end
			3942: begin
				if(in == 0) begin
					state<=5222;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=1333;
					out<=0;
				end
				if(in == 3) begin
					state<=7154;
					out<=1;
				end
				if(in == 4) begin
					state<=3265;
					out<=2;
				end
			end
			3943: begin
				if(in == 0) begin
					state<=5223;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=1334;
					out<=5;
				end
				if(in == 3) begin
					state<=7155;
					out<=6;
				end
				if(in == 4) begin
					state<=3266;
					out<=7;
				end
			end
			3944: begin
				if(in == 0) begin
					state<=5224;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=1335;
					out<=10;
				end
				if(in == 3) begin
					state<=7156;
					out<=11;
				end
				if(in == 4) begin
					state<=3267;
					out<=12;
				end
			end
			3945: begin
				if(in == 0) begin
					state<=5225;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=1336;
					out<=15;
				end
				if(in == 3) begin
					state<=7157;
					out<=16;
				end
				if(in == 4) begin
					state<=3268;
					out<=17;
				end
			end
			3946: begin
				if(in == 0) begin
					state<=5226;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=1337;
					out<=20;
				end
				if(in == 3) begin
					state<=7158;
					out<=21;
				end
				if(in == 4) begin
					state<=3269;
					out<=22;
				end
			end
			3947: begin
				if(in == 0) begin
					state<=5227;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=1338;
					out<=25;
				end
				if(in == 3) begin
					state<=7159;
					out<=26;
				end
				if(in == 4) begin
					state<=3270;
					out<=27;
				end
			end
			3948: begin
				if(in == 0) begin
					state<=5218;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=1329;
					out<=30;
				end
				if(in == 3) begin
					state<=7150;
					out<=31;
				end
				if(in == 4) begin
					state<=3261;
					out<=32;
				end
			end
			3949: begin
				if(in == 0) begin
					state<=3960;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=62;
					out<=35;
				end
				if(in == 3) begin
					state<=5949;
					out<=36;
				end
				if(in == 4) begin
					state<=2060;
					out<=37;
				end
			end
			3950: begin
				if(in == 0) begin
					state<=3961;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=63;
					out<=40;
				end
				if(in == 3) begin
					state<=5950;
					out<=41;
				end
				if(in == 4) begin
					state<=2061;
					out<=42;
				end
			end
			3951: begin
				if(in == 0) begin
					state<=3962;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=64;
					out<=45;
				end
				if(in == 3) begin
					state<=5951;
					out<=46;
				end
				if(in == 4) begin
					state<=2062;
					out<=47;
				end
			end
			3952: begin
				if(in == 0) begin
					state<=3963;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=65;
					out<=50;
				end
				if(in == 3) begin
					state<=5952;
					out<=51;
				end
				if(in == 4) begin
					state<=2063;
					out<=52;
				end
			end
			3953: begin
				if(in == 0) begin
					state<=3964;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=66;
					out<=55;
				end
				if(in == 3) begin
					state<=5953;
					out<=56;
				end
				if(in == 4) begin
					state<=2064;
					out<=57;
				end
			end
			3954: begin
				if(in == 0) begin
					state<=3965;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=67;
					out<=60;
				end
				if(in == 3) begin
					state<=5954;
					out<=61;
				end
				if(in == 4) begin
					state<=2065;
					out<=62;
				end
			end
			3955: begin
				if(in == 0) begin
					state<=3966;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=68;
					out<=65;
				end
				if(in == 3) begin
					state<=5955;
					out<=66;
				end
				if(in == 4) begin
					state<=2066;
					out<=67;
				end
			end
			3956: begin
				if(in == 0) begin
					state<=3967;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=69;
					out<=70;
				end
				if(in == 3) begin
					state<=5956;
					out<=71;
				end
				if(in == 4) begin
					state<=2067;
					out<=72;
				end
			end
			3957: begin
				if(in == 0) begin
					state<=3958;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=60;
					out<=75;
				end
				if(in == 3) begin
					state<=5947;
					out<=76;
				end
				if(in == 4) begin
					state<=2058;
					out<=77;
				end
			end
			3958: begin
				if(in == 0) begin
					state<=3969;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=71;
					out<=80;
				end
				if(in == 3) begin
					state<=5958;
					out<=81;
				end
				if(in == 4) begin
					state<=2069;
					out<=82;
				end
			end
			3959: begin
				if(in == 0) begin
					state<=3970;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=72;
					out<=85;
				end
				if(in == 3) begin
					state<=5959;
					out<=86;
				end
				if(in == 4) begin
					state<=2070;
					out<=87;
				end
			end
			3960: begin
				if(in == 0) begin
					state<=3971;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=73;
					out<=90;
				end
				if(in == 3) begin
					state<=5960;
					out<=91;
				end
				if(in == 4) begin
					state<=2071;
					out<=92;
				end
			end
			3961: begin
				if(in == 0) begin
					state<=3972;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=74;
					out<=95;
				end
				if(in == 3) begin
					state<=5961;
					out<=96;
				end
				if(in == 4) begin
					state<=2072;
					out<=97;
				end
			end
			3962: begin
				if(in == 0) begin
					state<=3973;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=75;
					out<=100;
				end
				if(in == 3) begin
					state<=5962;
					out<=101;
				end
				if(in == 4) begin
					state<=2073;
					out<=102;
				end
			end
			3963: begin
				if(in == 0) begin
					state<=3974;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=76;
					out<=105;
				end
				if(in == 3) begin
					state<=5963;
					out<=106;
				end
				if(in == 4) begin
					state<=2074;
					out<=107;
				end
			end
			3964: begin
				if(in == 0) begin
					state<=3975;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=77;
					out<=110;
				end
				if(in == 3) begin
					state<=5964;
					out<=111;
				end
				if(in == 4) begin
					state<=2075;
					out<=112;
				end
			end
			3965: begin
				if(in == 0) begin
					state<=3976;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=78;
					out<=115;
				end
				if(in == 3) begin
					state<=5965;
					out<=116;
				end
				if(in == 4) begin
					state<=2076;
					out<=117;
				end
			end
			3966: begin
				if(in == 0) begin
					state<=3977;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=79;
					out<=120;
				end
				if(in == 3) begin
					state<=5966;
					out<=121;
				end
				if(in == 4) begin
					state<=2077;
					out<=122;
				end
			end
			3967: begin
				if(in == 0) begin
					state<=3968;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=70;
					out<=125;
				end
				if(in == 3) begin
					state<=5957;
					out<=126;
				end
				if(in == 4) begin
					state<=2068;
					out<=127;
				end
			end
			3968: begin
				if(in == 0) begin
					state<=3979;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=81;
					out<=130;
				end
				if(in == 3) begin
					state<=5968;
					out<=131;
				end
				if(in == 4) begin
					state<=2079;
					out<=132;
				end
			end
			3969: begin
				if(in == 0) begin
					state<=3980;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=82;
					out<=135;
				end
				if(in == 3) begin
					state<=5969;
					out<=136;
				end
				if(in == 4) begin
					state<=2080;
					out<=137;
				end
			end
			3970: begin
				if(in == 0) begin
					state<=3981;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=83;
					out<=140;
				end
				if(in == 3) begin
					state<=5970;
					out<=141;
				end
				if(in == 4) begin
					state<=2081;
					out<=142;
				end
			end
			3971: begin
				if(in == 0) begin
					state<=3982;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=84;
					out<=145;
				end
				if(in == 3) begin
					state<=5971;
					out<=146;
				end
				if(in == 4) begin
					state<=2082;
					out<=147;
				end
			end
			3972: begin
				if(in == 0) begin
					state<=3983;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=85;
					out<=150;
				end
				if(in == 3) begin
					state<=5972;
					out<=151;
				end
				if(in == 4) begin
					state<=2083;
					out<=152;
				end
			end
			3973: begin
				if(in == 0) begin
					state<=3984;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=86;
					out<=155;
				end
				if(in == 3) begin
					state<=5973;
					out<=156;
				end
				if(in == 4) begin
					state<=2084;
					out<=157;
				end
			end
			3974: begin
				if(in == 0) begin
					state<=3985;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=87;
					out<=160;
				end
				if(in == 3) begin
					state<=5974;
					out<=161;
				end
				if(in == 4) begin
					state<=2085;
					out<=162;
				end
			end
			3975: begin
				if(in == 0) begin
					state<=3986;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=88;
					out<=165;
				end
				if(in == 3) begin
					state<=5975;
					out<=166;
				end
				if(in == 4) begin
					state<=2086;
					out<=167;
				end
			end
			3976: begin
				if(in == 0) begin
					state<=3987;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=89;
					out<=170;
				end
				if(in == 3) begin
					state<=5976;
					out<=171;
				end
				if(in == 4) begin
					state<=2087;
					out<=172;
				end
			end
			3977: begin
				if(in == 0) begin
					state<=3978;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=80;
					out<=175;
				end
				if(in == 3) begin
					state<=5967;
					out<=176;
				end
				if(in == 4) begin
					state<=2078;
					out<=177;
				end
			end
			3978: begin
				if(in == 0) begin
					state<=3989;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=91;
					out<=180;
				end
				if(in == 3) begin
					state<=5978;
					out<=181;
				end
				if(in == 4) begin
					state<=2089;
					out<=182;
				end
			end
			3979: begin
				if(in == 0) begin
					state<=3990;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=92;
					out<=185;
				end
				if(in == 3) begin
					state<=5979;
					out<=186;
				end
				if(in == 4) begin
					state<=2090;
					out<=187;
				end
			end
			3980: begin
				if(in == 0) begin
					state<=3991;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=93;
					out<=190;
				end
				if(in == 3) begin
					state<=5980;
					out<=191;
				end
				if(in == 4) begin
					state<=2091;
					out<=192;
				end
			end
			3981: begin
				if(in == 0) begin
					state<=3992;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=94;
					out<=195;
				end
				if(in == 3) begin
					state<=5981;
					out<=196;
				end
				if(in == 4) begin
					state<=2092;
					out<=197;
				end
			end
			3982: begin
				if(in == 0) begin
					state<=3993;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=95;
					out<=200;
				end
				if(in == 3) begin
					state<=5982;
					out<=201;
				end
				if(in == 4) begin
					state<=2093;
					out<=202;
				end
			end
			3983: begin
				if(in == 0) begin
					state<=3994;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=96;
					out<=205;
				end
				if(in == 3) begin
					state<=5983;
					out<=206;
				end
				if(in == 4) begin
					state<=2094;
					out<=207;
				end
			end
			3984: begin
				if(in == 0) begin
					state<=3995;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=97;
					out<=210;
				end
				if(in == 3) begin
					state<=5984;
					out<=211;
				end
				if(in == 4) begin
					state<=2095;
					out<=212;
				end
			end
			3985: begin
				if(in == 0) begin
					state<=3996;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=98;
					out<=215;
				end
				if(in == 3) begin
					state<=5985;
					out<=216;
				end
				if(in == 4) begin
					state<=2096;
					out<=217;
				end
			end
			3986: begin
				if(in == 0) begin
					state<=3997;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=99;
					out<=220;
				end
				if(in == 3) begin
					state<=5986;
					out<=221;
				end
				if(in == 4) begin
					state<=2097;
					out<=222;
				end
			end
			3987: begin
				if(in == 0) begin
					state<=3988;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=90;
					out<=225;
				end
				if(in == 3) begin
					state<=5977;
					out<=226;
				end
				if(in == 4) begin
					state<=2088;
					out<=227;
				end
			end
			3988: begin
				if(in == 0) begin
					state<=3999;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=101;
					out<=230;
				end
				if(in == 3) begin
					state<=5988;
					out<=231;
				end
				if(in == 4) begin
					state<=2099;
					out<=232;
				end
			end
			3989: begin
				if(in == 0) begin
					state<=4000;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=102;
					out<=235;
				end
				if(in == 3) begin
					state<=5989;
					out<=236;
				end
				if(in == 4) begin
					state<=2100;
					out<=237;
				end
			end
			3990: begin
				if(in == 0) begin
					state<=4001;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=103;
					out<=240;
				end
				if(in == 3) begin
					state<=5990;
					out<=241;
				end
				if(in == 4) begin
					state<=2101;
					out<=242;
				end
			end
			3991: begin
				if(in == 0) begin
					state<=4002;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=104;
					out<=245;
				end
				if(in == 3) begin
					state<=5991;
					out<=246;
				end
				if(in == 4) begin
					state<=2102;
					out<=247;
				end
			end
			3992: begin
				if(in == 0) begin
					state<=4003;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=105;
					out<=250;
				end
				if(in == 3) begin
					state<=5992;
					out<=251;
				end
				if(in == 4) begin
					state<=2103;
					out<=252;
				end
			end
			3993: begin
				if(in == 0) begin
					state<=4004;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=106;
					out<=255;
				end
				if(in == 3) begin
					state<=5993;
					out<=0;
				end
				if(in == 4) begin
					state<=2104;
					out<=1;
				end
			end
			3994: begin
				if(in == 0) begin
					state<=4005;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=107;
					out<=4;
				end
				if(in == 3) begin
					state<=5994;
					out<=5;
				end
				if(in == 4) begin
					state<=2105;
					out<=6;
				end
			end
			3995: begin
				if(in == 0) begin
					state<=4006;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=108;
					out<=9;
				end
				if(in == 3) begin
					state<=5995;
					out<=10;
				end
				if(in == 4) begin
					state<=2106;
					out<=11;
				end
			end
			3996: begin
				if(in == 0) begin
					state<=4007;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=109;
					out<=14;
				end
				if(in == 3) begin
					state<=5996;
					out<=15;
				end
				if(in == 4) begin
					state<=2107;
					out<=16;
				end
			end
			3997: begin
				if(in == 0) begin
					state<=3998;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=100;
					out<=19;
				end
				if(in == 3) begin
					state<=5987;
					out<=20;
				end
				if(in == 4) begin
					state<=2098;
					out<=21;
				end
			end
			3998: begin
				if(in == 0) begin
					state<=4009;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=111;
					out<=24;
				end
				if(in == 3) begin
					state<=5998;
					out<=25;
				end
				if(in == 4) begin
					state<=2109;
					out<=26;
				end
			end
			3999: begin
				if(in == 0) begin
					state<=4010;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=112;
					out<=29;
				end
				if(in == 3) begin
					state<=5999;
					out<=30;
				end
				if(in == 4) begin
					state<=2110;
					out<=31;
				end
			end
			4000: begin
				if(in == 0) begin
					state<=4011;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=113;
					out<=34;
				end
				if(in == 3) begin
					state<=6000;
					out<=35;
				end
				if(in == 4) begin
					state<=2111;
					out<=36;
				end
			end
			4001: begin
				if(in == 0) begin
					state<=4012;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=114;
					out<=39;
				end
				if(in == 3) begin
					state<=6001;
					out<=40;
				end
				if(in == 4) begin
					state<=2112;
					out<=41;
				end
			end
			4002: begin
				if(in == 0) begin
					state<=4013;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=115;
					out<=44;
				end
				if(in == 3) begin
					state<=6002;
					out<=45;
				end
				if(in == 4) begin
					state<=2113;
					out<=46;
				end
			end
			4003: begin
				if(in == 0) begin
					state<=4014;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=116;
					out<=49;
				end
				if(in == 3) begin
					state<=6003;
					out<=50;
				end
				if(in == 4) begin
					state<=2114;
					out<=51;
				end
			end
			4004: begin
				if(in == 0) begin
					state<=4015;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=117;
					out<=54;
				end
				if(in == 3) begin
					state<=6004;
					out<=55;
				end
				if(in == 4) begin
					state<=2115;
					out<=56;
				end
			end
			4005: begin
				if(in == 0) begin
					state<=4016;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=118;
					out<=59;
				end
				if(in == 3) begin
					state<=6005;
					out<=60;
				end
				if(in == 4) begin
					state<=2116;
					out<=61;
				end
			end
			4006: begin
				if(in == 0) begin
					state<=4017;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=119;
					out<=64;
				end
				if(in == 3) begin
					state<=6006;
					out<=65;
				end
				if(in == 4) begin
					state<=2117;
					out<=66;
				end
			end
			4007: begin
				if(in == 0) begin
					state<=4008;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=110;
					out<=69;
				end
				if(in == 3) begin
					state<=5997;
					out<=70;
				end
				if(in == 4) begin
					state<=2108;
					out<=71;
				end
			end
			4008: begin
				if(in == 0) begin
					state<=5250;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=1361;
					out<=74;
				end
				if(in == 3) begin
					state<=7182;
					out<=75;
				end
				if(in == 4) begin
					state<=3293;
					out<=76;
				end
			end
			4009: begin
				if(in == 0) begin
					state<=5251;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=1362;
					out<=79;
				end
				if(in == 3) begin
					state<=7183;
					out<=80;
				end
				if(in == 4) begin
					state<=3294;
					out<=81;
				end
			end
			4010: begin
				if(in == 0) begin
					state<=5252;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=1363;
					out<=84;
				end
				if(in == 3) begin
					state<=7184;
					out<=85;
				end
				if(in == 4) begin
					state<=3295;
					out<=86;
				end
			end
			4011: begin
				if(in == 0) begin
					state<=5253;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=1364;
					out<=89;
				end
				if(in == 3) begin
					state<=7185;
					out<=90;
				end
				if(in == 4) begin
					state<=3296;
					out<=91;
				end
			end
			4012: begin
				if(in == 0) begin
					state<=5254;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=1365;
					out<=94;
				end
				if(in == 3) begin
					state<=7186;
					out<=95;
				end
				if(in == 4) begin
					state<=3297;
					out<=96;
				end
			end
			4013: begin
				if(in == 0) begin
					state<=5255;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=1366;
					out<=99;
				end
				if(in == 3) begin
					state<=7187;
					out<=100;
				end
				if(in == 4) begin
					state<=3298;
					out<=101;
				end
			end
			4014: begin
				if(in == 0) begin
					state<=5256;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=1367;
					out<=104;
				end
				if(in == 3) begin
					state<=7188;
					out<=105;
				end
				if(in == 4) begin
					state<=3299;
					out<=106;
				end
			end
			4015: begin
				if(in == 0) begin
					state<=5257;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=1368;
					out<=109;
				end
				if(in == 3) begin
					state<=7189;
					out<=110;
				end
				if(in == 4) begin
					state<=3300;
					out<=111;
				end
			end
			4016: begin
				if(in == 0) begin
					state<=5258;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=1369;
					out<=114;
				end
				if(in == 3) begin
					state<=7190;
					out<=115;
				end
				if(in == 4) begin
					state<=3301;
					out<=116;
				end
			end
			4017: begin
				if(in == 0) begin
					state<=5249;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=1360;
					out<=119;
				end
				if(in == 3) begin
					state<=7181;
					out<=120;
				end
				if(in == 4) begin
					state<=3292;
					out<=121;
				end
			end
			4018: begin
				if(in == 0) begin
					state<=4029;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=131;
					out<=124;
				end
				if(in == 3) begin
					state<=6018;
					out<=125;
				end
				if(in == 4) begin
					state<=2129;
					out<=126;
				end
			end
			4019: begin
				if(in == 0) begin
					state<=4030;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=132;
					out<=129;
				end
				if(in == 3) begin
					state<=6019;
					out<=130;
				end
				if(in == 4) begin
					state<=2130;
					out<=131;
				end
			end
			4020: begin
				if(in == 0) begin
					state<=4031;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=133;
					out<=134;
				end
				if(in == 3) begin
					state<=6020;
					out<=135;
				end
				if(in == 4) begin
					state<=2131;
					out<=136;
				end
			end
			4021: begin
				if(in == 0) begin
					state<=4032;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=134;
					out<=139;
				end
				if(in == 3) begin
					state<=6021;
					out<=140;
				end
				if(in == 4) begin
					state<=2132;
					out<=141;
				end
			end
			4022: begin
				if(in == 0) begin
					state<=4033;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=135;
					out<=144;
				end
				if(in == 3) begin
					state<=6022;
					out<=145;
				end
				if(in == 4) begin
					state<=2133;
					out<=146;
				end
			end
			4023: begin
				if(in == 0) begin
					state<=4034;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=136;
					out<=149;
				end
				if(in == 3) begin
					state<=6023;
					out<=150;
				end
				if(in == 4) begin
					state<=2134;
					out<=151;
				end
			end
			4024: begin
				if(in == 0) begin
					state<=4035;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=137;
					out<=154;
				end
				if(in == 3) begin
					state<=6024;
					out<=155;
				end
				if(in == 4) begin
					state<=2135;
					out<=156;
				end
			end
			4025: begin
				if(in == 0) begin
					state<=4036;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=138;
					out<=159;
				end
				if(in == 3) begin
					state<=6025;
					out<=160;
				end
				if(in == 4) begin
					state<=2136;
					out<=161;
				end
			end
			4026: begin
				if(in == 0) begin
					state<=4027;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=129;
					out<=164;
				end
				if(in == 3) begin
					state<=6016;
					out<=165;
				end
				if(in == 4) begin
					state<=2127;
					out<=166;
				end
			end
			4027: begin
				if(in == 0) begin
					state<=4038;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=140;
					out<=169;
				end
				if(in == 3) begin
					state<=6027;
					out<=170;
				end
				if(in == 4) begin
					state<=2138;
					out<=171;
				end
			end
			4028: begin
				if(in == 0) begin
					state<=4039;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=141;
					out<=174;
				end
				if(in == 3) begin
					state<=6028;
					out<=175;
				end
				if(in == 4) begin
					state<=2139;
					out<=176;
				end
			end
			4029: begin
				if(in == 0) begin
					state<=4040;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=142;
					out<=179;
				end
				if(in == 3) begin
					state<=6029;
					out<=180;
				end
				if(in == 4) begin
					state<=2140;
					out<=181;
				end
			end
			4030: begin
				if(in == 0) begin
					state<=4041;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=143;
					out<=184;
				end
				if(in == 3) begin
					state<=6030;
					out<=185;
				end
				if(in == 4) begin
					state<=2141;
					out<=186;
				end
			end
			4031: begin
				if(in == 0) begin
					state<=4042;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=144;
					out<=189;
				end
				if(in == 3) begin
					state<=6031;
					out<=190;
				end
				if(in == 4) begin
					state<=2142;
					out<=191;
				end
			end
			4032: begin
				if(in == 0) begin
					state<=4043;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=145;
					out<=194;
				end
				if(in == 3) begin
					state<=6032;
					out<=195;
				end
				if(in == 4) begin
					state<=2143;
					out<=196;
				end
			end
			4033: begin
				if(in == 0) begin
					state<=4044;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=146;
					out<=199;
				end
				if(in == 3) begin
					state<=6033;
					out<=200;
				end
				if(in == 4) begin
					state<=2144;
					out<=201;
				end
			end
			4034: begin
				if(in == 0) begin
					state<=4045;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=147;
					out<=204;
				end
				if(in == 3) begin
					state<=6034;
					out<=205;
				end
				if(in == 4) begin
					state<=2145;
					out<=206;
				end
			end
			4035: begin
				if(in == 0) begin
					state<=4046;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=148;
					out<=209;
				end
				if(in == 3) begin
					state<=6035;
					out<=210;
				end
				if(in == 4) begin
					state<=2146;
					out<=211;
				end
			end
			4036: begin
				if(in == 0) begin
					state<=4037;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=139;
					out<=214;
				end
				if(in == 3) begin
					state<=6026;
					out<=215;
				end
				if(in == 4) begin
					state<=2137;
					out<=216;
				end
			end
			4037: begin
				if(in == 0) begin
					state<=4048;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=150;
					out<=219;
				end
				if(in == 3) begin
					state<=6037;
					out<=220;
				end
				if(in == 4) begin
					state<=2148;
					out<=221;
				end
			end
			4038: begin
				if(in == 0) begin
					state<=4049;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=151;
					out<=224;
				end
				if(in == 3) begin
					state<=6038;
					out<=225;
				end
				if(in == 4) begin
					state<=2149;
					out<=226;
				end
			end
			4039: begin
				if(in == 0) begin
					state<=4050;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=152;
					out<=229;
				end
				if(in == 3) begin
					state<=6039;
					out<=230;
				end
				if(in == 4) begin
					state<=2150;
					out<=231;
				end
			end
			4040: begin
				if(in == 0) begin
					state<=4051;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=153;
					out<=234;
				end
				if(in == 3) begin
					state<=6040;
					out<=235;
				end
				if(in == 4) begin
					state<=2151;
					out<=236;
				end
			end
			4041: begin
				if(in == 0) begin
					state<=4052;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=154;
					out<=239;
				end
				if(in == 3) begin
					state<=6041;
					out<=240;
				end
				if(in == 4) begin
					state<=2152;
					out<=241;
				end
			end
			4042: begin
				if(in == 0) begin
					state<=4053;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=155;
					out<=244;
				end
				if(in == 3) begin
					state<=6042;
					out<=245;
				end
				if(in == 4) begin
					state<=2153;
					out<=246;
				end
			end
			4043: begin
				if(in == 0) begin
					state<=4054;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=156;
					out<=249;
				end
				if(in == 3) begin
					state<=6043;
					out<=250;
				end
				if(in == 4) begin
					state<=2154;
					out<=251;
				end
			end
			4044: begin
				if(in == 0) begin
					state<=4055;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=157;
					out<=254;
				end
				if(in == 3) begin
					state<=6044;
					out<=255;
				end
				if(in == 4) begin
					state<=2155;
					out<=0;
				end
			end
			4045: begin
				if(in == 0) begin
					state<=4056;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=158;
					out<=3;
				end
				if(in == 3) begin
					state<=6045;
					out<=4;
				end
				if(in == 4) begin
					state<=2156;
					out<=5;
				end
			end
			4046: begin
				if(in == 0) begin
					state<=4047;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=149;
					out<=8;
				end
				if(in == 3) begin
					state<=6036;
					out<=9;
				end
				if(in == 4) begin
					state<=2147;
					out<=10;
				end
			end
			4047: begin
				if(in == 0) begin
					state<=4058;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=160;
					out<=13;
				end
				if(in == 3) begin
					state<=6047;
					out<=14;
				end
				if(in == 4) begin
					state<=2158;
					out<=15;
				end
			end
			4048: begin
				if(in == 0) begin
					state<=4059;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=161;
					out<=18;
				end
				if(in == 3) begin
					state<=6048;
					out<=19;
				end
				if(in == 4) begin
					state<=2159;
					out<=20;
				end
			end
			4049: begin
				if(in == 0) begin
					state<=4060;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=162;
					out<=23;
				end
				if(in == 3) begin
					state<=6049;
					out<=24;
				end
				if(in == 4) begin
					state<=2160;
					out<=25;
				end
			end
			4050: begin
				if(in == 0) begin
					state<=4061;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=163;
					out<=28;
				end
				if(in == 3) begin
					state<=6050;
					out<=29;
				end
				if(in == 4) begin
					state<=2161;
					out<=30;
				end
			end
			4051: begin
				if(in == 0) begin
					state<=4062;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=164;
					out<=33;
				end
				if(in == 3) begin
					state<=6051;
					out<=34;
				end
				if(in == 4) begin
					state<=2162;
					out<=35;
				end
			end
			4052: begin
				if(in == 0) begin
					state<=4063;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=165;
					out<=38;
				end
				if(in == 3) begin
					state<=6052;
					out<=39;
				end
				if(in == 4) begin
					state<=2163;
					out<=40;
				end
			end
			4053: begin
				if(in == 0) begin
					state<=4064;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=166;
					out<=43;
				end
				if(in == 3) begin
					state<=6053;
					out<=44;
				end
				if(in == 4) begin
					state<=2164;
					out<=45;
				end
			end
			4054: begin
				if(in == 0) begin
					state<=4065;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=167;
					out<=48;
				end
				if(in == 3) begin
					state<=6054;
					out<=49;
				end
				if(in == 4) begin
					state<=2165;
					out<=50;
				end
			end
			4055: begin
				if(in == 0) begin
					state<=4066;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=168;
					out<=53;
				end
				if(in == 3) begin
					state<=6055;
					out<=54;
				end
				if(in == 4) begin
					state<=2166;
					out<=55;
				end
			end
			4056: begin
				if(in == 0) begin
					state<=4057;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=159;
					out<=58;
				end
				if(in == 3) begin
					state<=6046;
					out<=59;
				end
				if(in == 4) begin
					state<=2157;
					out<=60;
				end
			end
			4057: begin
				if(in == 0) begin
					state<=4068;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=170;
					out<=63;
				end
				if(in == 3) begin
					state<=6057;
					out<=64;
				end
				if(in == 4) begin
					state<=2168;
					out<=65;
				end
			end
			4058: begin
				if(in == 0) begin
					state<=4069;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=171;
					out<=68;
				end
				if(in == 3) begin
					state<=6058;
					out<=69;
				end
				if(in == 4) begin
					state<=2169;
					out<=70;
				end
			end
			4059: begin
				if(in == 0) begin
					state<=4070;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=172;
					out<=73;
				end
				if(in == 3) begin
					state<=6059;
					out<=74;
				end
				if(in == 4) begin
					state<=2170;
					out<=75;
				end
			end
			4060: begin
				if(in == 0) begin
					state<=4071;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=173;
					out<=78;
				end
				if(in == 3) begin
					state<=6060;
					out<=79;
				end
				if(in == 4) begin
					state<=2171;
					out<=80;
				end
			end
			4061: begin
				if(in == 0) begin
					state<=4072;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=174;
					out<=83;
				end
				if(in == 3) begin
					state<=6061;
					out<=84;
				end
				if(in == 4) begin
					state<=2172;
					out<=85;
				end
			end
			4062: begin
				if(in == 0) begin
					state<=4073;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=175;
					out<=88;
				end
				if(in == 3) begin
					state<=6062;
					out<=89;
				end
				if(in == 4) begin
					state<=2173;
					out<=90;
				end
			end
			4063: begin
				if(in == 0) begin
					state<=4074;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=176;
					out<=93;
				end
				if(in == 3) begin
					state<=6063;
					out<=94;
				end
				if(in == 4) begin
					state<=2174;
					out<=95;
				end
			end
			4064: begin
				if(in == 0) begin
					state<=4075;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=177;
					out<=98;
				end
				if(in == 3) begin
					state<=6064;
					out<=99;
				end
				if(in == 4) begin
					state<=2175;
					out<=100;
				end
			end
			4065: begin
				if(in == 0) begin
					state<=4076;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=178;
					out<=103;
				end
				if(in == 3) begin
					state<=6065;
					out<=104;
				end
				if(in == 4) begin
					state<=2176;
					out<=105;
				end
			end
			4066: begin
				if(in == 0) begin
					state<=4067;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=169;
					out<=108;
				end
				if(in == 3) begin
					state<=6056;
					out<=109;
				end
				if(in == 4) begin
					state<=2167;
					out<=110;
				end
			end
			4067: begin
				if(in == 0) begin
					state<=4078;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=180;
					out<=113;
				end
				if(in == 3) begin
					state<=6067;
					out<=114;
				end
				if(in == 4) begin
					state<=2178;
					out<=115;
				end
			end
			4068: begin
				if(in == 0) begin
					state<=4079;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=181;
					out<=118;
				end
				if(in == 3) begin
					state<=6068;
					out<=119;
				end
				if(in == 4) begin
					state<=2179;
					out<=120;
				end
			end
			4069: begin
				if(in == 0) begin
					state<=4080;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=182;
					out<=123;
				end
				if(in == 3) begin
					state<=6069;
					out<=124;
				end
				if(in == 4) begin
					state<=2180;
					out<=125;
				end
			end
			4070: begin
				if(in == 0) begin
					state<=4081;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=183;
					out<=128;
				end
				if(in == 3) begin
					state<=6070;
					out<=129;
				end
				if(in == 4) begin
					state<=2181;
					out<=130;
				end
			end
			4071: begin
				if(in == 0) begin
					state<=4082;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=184;
					out<=133;
				end
				if(in == 3) begin
					state<=6071;
					out<=134;
				end
				if(in == 4) begin
					state<=2182;
					out<=135;
				end
			end
			4072: begin
				if(in == 0) begin
					state<=4083;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=185;
					out<=138;
				end
				if(in == 3) begin
					state<=6072;
					out<=139;
				end
				if(in == 4) begin
					state<=2183;
					out<=140;
				end
			end
			4073: begin
				if(in == 0) begin
					state<=4084;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=186;
					out<=143;
				end
				if(in == 3) begin
					state<=6073;
					out<=144;
				end
				if(in == 4) begin
					state<=2184;
					out<=145;
				end
			end
			4074: begin
				if(in == 0) begin
					state<=4085;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=187;
					out<=148;
				end
				if(in == 3) begin
					state<=6074;
					out<=149;
				end
				if(in == 4) begin
					state<=2185;
					out<=150;
				end
			end
			4075: begin
				if(in == 0) begin
					state<=4086;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=188;
					out<=153;
				end
				if(in == 3) begin
					state<=6075;
					out<=154;
				end
				if(in == 4) begin
					state<=2186;
					out<=155;
				end
			end
			4076: begin
				if(in == 0) begin
					state<=4077;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=179;
					out<=158;
				end
				if(in == 3) begin
					state<=6066;
					out<=159;
				end
				if(in == 4) begin
					state<=2177;
					out<=160;
				end
			end
			4077: begin
				if(in == 0) begin
					state<=5281;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=1392;
					out<=163;
				end
				if(in == 3) begin
					state<=7213;
					out<=164;
				end
				if(in == 4) begin
					state<=3324;
					out<=165;
				end
			end
			4078: begin
				if(in == 0) begin
					state<=5282;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=1393;
					out<=168;
				end
				if(in == 3) begin
					state<=7214;
					out<=169;
				end
				if(in == 4) begin
					state<=3325;
					out<=170;
				end
			end
			4079: begin
				if(in == 0) begin
					state<=5283;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=1394;
					out<=173;
				end
				if(in == 3) begin
					state<=7215;
					out<=174;
				end
				if(in == 4) begin
					state<=3326;
					out<=175;
				end
			end
			4080: begin
				if(in == 0) begin
					state<=5284;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=1395;
					out<=178;
				end
				if(in == 3) begin
					state<=7216;
					out<=179;
				end
				if(in == 4) begin
					state<=3327;
					out<=180;
				end
			end
			4081: begin
				if(in == 0) begin
					state<=5285;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=1396;
					out<=183;
				end
				if(in == 3) begin
					state<=7217;
					out<=184;
				end
				if(in == 4) begin
					state<=3328;
					out<=185;
				end
			end
			4082: begin
				if(in == 0) begin
					state<=5286;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=1397;
					out<=188;
				end
				if(in == 3) begin
					state<=7218;
					out<=189;
				end
				if(in == 4) begin
					state<=3329;
					out<=190;
				end
			end
			4083: begin
				if(in == 0) begin
					state<=5287;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=1398;
					out<=193;
				end
				if(in == 3) begin
					state<=7219;
					out<=194;
				end
				if(in == 4) begin
					state<=3330;
					out<=195;
				end
			end
			4084: begin
				if(in == 0) begin
					state<=5288;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=1399;
					out<=198;
				end
				if(in == 3) begin
					state<=7220;
					out<=199;
				end
				if(in == 4) begin
					state<=3331;
					out<=200;
				end
			end
			4085: begin
				if(in == 0) begin
					state<=5289;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=1400;
					out<=203;
				end
				if(in == 3) begin
					state<=7221;
					out<=204;
				end
				if(in == 4) begin
					state<=3332;
					out<=205;
				end
			end
			4086: begin
				if(in == 0) begin
					state<=5280;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=1391;
					out<=208;
				end
				if(in == 3) begin
					state<=7212;
					out<=209;
				end
				if(in == 4) begin
					state<=3323;
					out<=210;
				end
			end
			4087: begin
				if(in == 0) begin
					state<=4098;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=200;
					out<=213;
				end
				if(in == 3) begin
					state<=6087;
					out<=214;
				end
				if(in == 4) begin
					state<=2198;
					out<=215;
				end
			end
			4088: begin
				if(in == 0) begin
					state<=4099;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=201;
					out<=218;
				end
				if(in == 3) begin
					state<=6088;
					out<=219;
				end
				if(in == 4) begin
					state<=2199;
					out<=220;
				end
			end
			4089: begin
				if(in == 0) begin
					state<=4100;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=202;
					out<=223;
				end
				if(in == 3) begin
					state<=6089;
					out<=224;
				end
				if(in == 4) begin
					state<=2200;
					out<=225;
				end
			end
			4090: begin
				if(in == 0) begin
					state<=4101;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=203;
					out<=228;
				end
				if(in == 3) begin
					state<=6090;
					out<=229;
				end
				if(in == 4) begin
					state<=2201;
					out<=230;
				end
			end
			4091: begin
				if(in == 0) begin
					state<=4102;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=204;
					out<=233;
				end
				if(in == 3) begin
					state<=6091;
					out<=234;
				end
				if(in == 4) begin
					state<=2202;
					out<=235;
				end
			end
			4092: begin
				if(in == 0) begin
					state<=4103;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=205;
					out<=238;
				end
				if(in == 3) begin
					state<=6092;
					out<=239;
				end
				if(in == 4) begin
					state<=2203;
					out<=240;
				end
			end
			4093: begin
				if(in == 0) begin
					state<=4104;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=206;
					out<=243;
				end
				if(in == 3) begin
					state<=6093;
					out<=244;
				end
				if(in == 4) begin
					state<=2204;
					out<=245;
				end
			end
			4094: begin
				if(in == 0) begin
					state<=4105;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=207;
					out<=248;
				end
				if(in == 3) begin
					state<=6094;
					out<=249;
				end
				if(in == 4) begin
					state<=2205;
					out<=250;
				end
			end
			4095: begin
				if(in == 0) begin
					state<=4096;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=198;
					out<=253;
				end
				if(in == 3) begin
					state<=6085;
					out<=254;
				end
				if(in == 4) begin
					state<=2196;
					out<=255;
				end
			end
			4096: begin
				if(in == 0) begin
					state<=4107;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=209;
					out<=2;
				end
				if(in == 3) begin
					state<=6096;
					out<=3;
				end
				if(in == 4) begin
					state<=2207;
					out<=4;
				end
			end
			4097: begin
				if(in == 0) begin
					state<=4108;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=210;
					out<=7;
				end
				if(in == 3) begin
					state<=6097;
					out<=8;
				end
				if(in == 4) begin
					state<=2208;
					out<=9;
				end
			end
			4098: begin
				if(in == 0) begin
					state<=4109;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=211;
					out<=12;
				end
				if(in == 3) begin
					state<=6098;
					out<=13;
				end
				if(in == 4) begin
					state<=2209;
					out<=14;
				end
			end
			4099: begin
				if(in == 0) begin
					state<=4110;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=212;
					out<=17;
				end
				if(in == 3) begin
					state<=6099;
					out<=18;
				end
				if(in == 4) begin
					state<=2210;
					out<=19;
				end
			end
			4100: begin
				if(in == 0) begin
					state<=4111;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=213;
					out<=22;
				end
				if(in == 3) begin
					state<=6100;
					out<=23;
				end
				if(in == 4) begin
					state<=2211;
					out<=24;
				end
			end
			4101: begin
				if(in == 0) begin
					state<=4112;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=214;
					out<=27;
				end
				if(in == 3) begin
					state<=6101;
					out<=28;
				end
				if(in == 4) begin
					state<=2212;
					out<=29;
				end
			end
			4102: begin
				if(in == 0) begin
					state<=4113;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=215;
					out<=32;
				end
				if(in == 3) begin
					state<=6102;
					out<=33;
				end
				if(in == 4) begin
					state<=2213;
					out<=34;
				end
			end
			4103: begin
				if(in == 0) begin
					state<=4114;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=216;
					out<=37;
				end
				if(in == 3) begin
					state<=6103;
					out<=38;
				end
				if(in == 4) begin
					state<=2214;
					out<=39;
				end
			end
			4104: begin
				if(in == 0) begin
					state<=4115;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=217;
					out<=42;
				end
				if(in == 3) begin
					state<=6104;
					out<=43;
				end
				if(in == 4) begin
					state<=2215;
					out<=44;
				end
			end
			4105: begin
				if(in == 0) begin
					state<=4106;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=208;
					out<=47;
				end
				if(in == 3) begin
					state<=6095;
					out<=48;
				end
				if(in == 4) begin
					state<=2206;
					out<=49;
				end
			end
			4106: begin
				if(in == 0) begin
					state<=4117;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=219;
					out<=52;
				end
				if(in == 3) begin
					state<=6106;
					out<=53;
				end
				if(in == 4) begin
					state<=2217;
					out<=54;
				end
			end
			4107: begin
				if(in == 0) begin
					state<=4118;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=220;
					out<=57;
				end
				if(in == 3) begin
					state<=6107;
					out<=58;
				end
				if(in == 4) begin
					state<=2218;
					out<=59;
				end
			end
			4108: begin
				if(in == 0) begin
					state<=4119;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=221;
					out<=62;
				end
				if(in == 3) begin
					state<=6108;
					out<=63;
				end
				if(in == 4) begin
					state<=2219;
					out<=64;
				end
			end
			4109: begin
				if(in == 0) begin
					state<=4120;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=222;
					out<=67;
				end
				if(in == 3) begin
					state<=6109;
					out<=68;
				end
				if(in == 4) begin
					state<=2220;
					out<=69;
				end
			end
			4110: begin
				if(in == 0) begin
					state<=4121;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=223;
					out<=72;
				end
				if(in == 3) begin
					state<=6110;
					out<=73;
				end
				if(in == 4) begin
					state<=2221;
					out<=74;
				end
			end
			4111: begin
				if(in == 0) begin
					state<=4122;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=224;
					out<=77;
				end
				if(in == 3) begin
					state<=6111;
					out<=78;
				end
				if(in == 4) begin
					state<=2222;
					out<=79;
				end
			end
			4112: begin
				if(in == 0) begin
					state<=4123;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=225;
					out<=82;
				end
				if(in == 3) begin
					state<=6112;
					out<=83;
				end
				if(in == 4) begin
					state<=2223;
					out<=84;
				end
			end
			4113: begin
				if(in == 0) begin
					state<=4124;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=226;
					out<=87;
				end
				if(in == 3) begin
					state<=6113;
					out<=88;
				end
				if(in == 4) begin
					state<=2224;
					out<=89;
				end
			end
			4114: begin
				if(in == 0) begin
					state<=4125;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=227;
					out<=92;
				end
				if(in == 3) begin
					state<=6114;
					out<=93;
				end
				if(in == 4) begin
					state<=2225;
					out<=94;
				end
			end
			4115: begin
				if(in == 0) begin
					state<=4116;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=218;
					out<=97;
				end
				if(in == 3) begin
					state<=6105;
					out<=98;
				end
				if(in == 4) begin
					state<=2216;
					out<=99;
				end
			end
			4116: begin
				if(in == 0) begin
					state<=4127;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=229;
					out<=102;
				end
				if(in == 3) begin
					state<=6116;
					out<=103;
				end
				if(in == 4) begin
					state<=2227;
					out<=104;
				end
			end
			4117: begin
				if(in == 0) begin
					state<=4128;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=230;
					out<=107;
				end
				if(in == 3) begin
					state<=6117;
					out<=108;
				end
				if(in == 4) begin
					state<=2228;
					out<=109;
				end
			end
			4118: begin
				if(in == 0) begin
					state<=4129;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=231;
					out<=112;
				end
				if(in == 3) begin
					state<=6118;
					out<=113;
				end
				if(in == 4) begin
					state<=2229;
					out<=114;
				end
			end
			4119: begin
				if(in == 0) begin
					state<=4130;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=232;
					out<=117;
				end
				if(in == 3) begin
					state<=6119;
					out<=118;
				end
				if(in == 4) begin
					state<=2230;
					out<=119;
				end
			end
			4120: begin
				if(in == 0) begin
					state<=4131;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=233;
					out<=122;
				end
				if(in == 3) begin
					state<=6120;
					out<=123;
				end
				if(in == 4) begin
					state<=2231;
					out<=124;
				end
			end
			4121: begin
				if(in == 0) begin
					state<=4132;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=234;
					out<=127;
				end
				if(in == 3) begin
					state<=6121;
					out<=128;
				end
				if(in == 4) begin
					state<=2232;
					out<=129;
				end
			end
			4122: begin
				if(in == 0) begin
					state<=4133;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=235;
					out<=132;
				end
				if(in == 3) begin
					state<=6122;
					out<=133;
				end
				if(in == 4) begin
					state<=2233;
					out<=134;
				end
			end
			4123: begin
				if(in == 0) begin
					state<=4134;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=236;
					out<=137;
				end
				if(in == 3) begin
					state<=6123;
					out<=138;
				end
				if(in == 4) begin
					state<=2234;
					out<=139;
				end
			end
			4124: begin
				if(in == 0) begin
					state<=4135;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=237;
					out<=142;
				end
				if(in == 3) begin
					state<=6124;
					out<=143;
				end
				if(in == 4) begin
					state<=2235;
					out<=144;
				end
			end
			4125: begin
				if(in == 0) begin
					state<=4126;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=228;
					out<=147;
				end
				if(in == 3) begin
					state<=6115;
					out<=148;
				end
				if(in == 4) begin
					state<=2226;
					out<=149;
				end
			end
			4126: begin
				if(in == 0) begin
					state<=4137;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=239;
					out<=152;
				end
				if(in == 3) begin
					state<=6126;
					out<=153;
				end
				if(in == 4) begin
					state<=2237;
					out<=154;
				end
			end
			4127: begin
				if(in == 0) begin
					state<=4138;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=240;
					out<=157;
				end
				if(in == 3) begin
					state<=6127;
					out<=158;
				end
				if(in == 4) begin
					state<=2238;
					out<=159;
				end
			end
			4128: begin
				if(in == 0) begin
					state<=4139;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=241;
					out<=162;
				end
				if(in == 3) begin
					state<=6128;
					out<=163;
				end
				if(in == 4) begin
					state<=2239;
					out<=164;
				end
			end
			4129: begin
				if(in == 0) begin
					state<=4140;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=242;
					out<=167;
				end
				if(in == 3) begin
					state<=6129;
					out<=168;
				end
				if(in == 4) begin
					state<=2240;
					out<=169;
				end
			end
			4130: begin
				if(in == 0) begin
					state<=4141;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=243;
					out<=172;
				end
				if(in == 3) begin
					state<=6130;
					out<=173;
				end
				if(in == 4) begin
					state<=2241;
					out<=174;
				end
			end
			4131: begin
				if(in == 0) begin
					state<=4142;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=244;
					out<=177;
				end
				if(in == 3) begin
					state<=6131;
					out<=178;
				end
				if(in == 4) begin
					state<=2242;
					out<=179;
				end
			end
			4132: begin
				if(in == 0) begin
					state<=4143;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=245;
					out<=182;
				end
				if(in == 3) begin
					state<=6132;
					out<=183;
				end
				if(in == 4) begin
					state<=2243;
					out<=184;
				end
			end
			4133: begin
				if(in == 0) begin
					state<=4144;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=246;
					out<=187;
				end
				if(in == 3) begin
					state<=6133;
					out<=188;
				end
				if(in == 4) begin
					state<=2244;
					out<=189;
				end
			end
			4134: begin
				if(in == 0) begin
					state<=4145;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=247;
					out<=192;
				end
				if(in == 3) begin
					state<=6134;
					out<=193;
				end
				if(in == 4) begin
					state<=2245;
					out<=194;
				end
			end
			4135: begin
				if(in == 0) begin
					state<=4136;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=238;
					out<=197;
				end
				if(in == 3) begin
					state<=6125;
					out<=198;
				end
				if(in == 4) begin
					state<=2236;
					out<=199;
				end
			end
			4136: begin
				if(in == 0) begin
					state<=4147;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=249;
					out<=202;
				end
				if(in == 3) begin
					state<=6136;
					out<=203;
				end
				if(in == 4) begin
					state<=2247;
					out<=204;
				end
			end
			4137: begin
				if(in == 0) begin
					state<=4148;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=250;
					out<=207;
				end
				if(in == 3) begin
					state<=6137;
					out<=208;
				end
				if(in == 4) begin
					state<=2248;
					out<=209;
				end
			end
			4138: begin
				if(in == 0) begin
					state<=4149;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=251;
					out<=212;
				end
				if(in == 3) begin
					state<=6138;
					out<=213;
				end
				if(in == 4) begin
					state<=2249;
					out<=214;
				end
			end
			4139: begin
				if(in == 0) begin
					state<=4150;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=252;
					out<=217;
				end
				if(in == 3) begin
					state<=6139;
					out<=218;
				end
				if(in == 4) begin
					state<=2250;
					out<=219;
				end
			end
			4140: begin
				if(in == 0) begin
					state<=4151;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=253;
					out<=222;
				end
				if(in == 3) begin
					state<=6140;
					out<=223;
				end
				if(in == 4) begin
					state<=2251;
					out<=224;
				end
			end
			4141: begin
				if(in == 0) begin
					state<=4152;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=254;
					out<=227;
				end
				if(in == 3) begin
					state<=6141;
					out<=228;
				end
				if(in == 4) begin
					state<=2252;
					out<=229;
				end
			end
			4142: begin
				if(in == 0) begin
					state<=4153;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=255;
					out<=232;
				end
				if(in == 3) begin
					state<=6142;
					out<=233;
				end
				if(in == 4) begin
					state<=2253;
					out<=234;
				end
			end
			4143: begin
				if(in == 0) begin
					state<=4154;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=256;
					out<=237;
				end
				if(in == 3) begin
					state<=6143;
					out<=238;
				end
				if(in == 4) begin
					state<=2254;
					out<=239;
				end
			end
			4144: begin
				if(in == 0) begin
					state<=4155;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=257;
					out<=242;
				end
				if(in == 3) begin
					state<=6144;
					out<=243;
				end
				if(in == 4) begin
					state<=2255;
					out<=244;
				end
			end
			4145: begin
				if(in == 0) begin
					state<=4146;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=248;
					out<=247;
				end
				if(in == 3) begin
					state<=6135;
					out<=248;
				end
				if(in == 4) begin
					state<=2246;
					out<=249;
				end
			end
			4146: begin
				if(in == 0) begin
					state<=5312;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=1423;
					out<=252;
				end
				if(in == 3) begin
					state<=7244;
					out<=253;
				end
				if(in == 4) begin
					state<=3355;
					out<=254;
				end
			end
			4147: begin
				if(in == 0) begin
					state<=5313;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=1424;
					out<=1;
				end
				if(in == 3) begin
					state<=7245;
					out<=2;
				end
				if(in == 4) begin
					state<=3356;
					out<=3;
				end
			end
			4148: begin
				if(in == 0) begin
					state<=5314;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=1425;
					out<=6;
				end
				if(in == 3) begin
					state<=7246;
					out<=7;
				end
				if(in == 4) begin
					state<=3357;
					out<=8;
				end
			end
			4149: begin
				if(in == 0) begin
					state<=5315;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=1426;
					out<=11;
				end
				if(in == 3) begin
					state<=7247;
					out<=12;
				end
				if(in == 4) begin
					state<=3358;
					out<=13;
				end
			end
			4150: begin
				if(in == 0) begin
					state<=5316;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=1427;
					out<=16;
				end
				if(in == 3) begin
					state<=7248;
					out<=17;
				end
				if(in == 4) begin
					state<=3359;
					out<=18;
				end
			end
			4151: begin
				if(in == 0) begin
					state<=5317;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=1428;
					out<=21;
				end
				if(in == 3) begin
					state<=7249;
					out<=22;
				end
				if(in == 4) begin
					state<=3360;
					out<=23;
				end
			end
			4152: begin
				if(in == 0) begin
					state<=5318;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=1429;
					out<=26;
				end
				if(in == 3) begin
					state<=7250;
					out<=27;
				end
				if(in == 4) begin
					state<=3361;
					out<=28;
				end
			end
			4153: begin
				if(in == 0) begin
					state<=5319;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=1430;
					out<=31;
				end
				if(in == 3) begin
					state<=7251;
					out<=32;
				end
				if(in == 4) begin
					state<=3362;
					out<=33;
				end
			end
			4154: begin
				if(in == 0) begin
					state<=5320;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=1431;
					out<=36;
				end
				if(in == 3) begin
					state<=7252;
					out<=37;
				end
				if(in == 4) begin
					state<=3363;
					out<=38;
				end
			end
			4155: begin
				if(in == 0) begin
					state<=5311;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=1422;
					out<=41;
				end
				if(in == 3) begin
					state<=7243;
					out<=42;
				end
				if(in == 4) begin
					state<=3354;
					out<=43;
				end
			end
			4156: begin
				if(in == 0) begin
					state<=4167;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=269;
					out<=46;
				end
				if(in == 3) begin
					state<=6156;
					out<=47;
				end
				if(in == 4) begin
					state<=2267;
					out<=48;
				end
			end
			4157: begin
				if(in == 0) begin
					state<=4168;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=270;
					out<=51;
				end
				if(in == 3) begin
					state<=6157;
					out<=52;
				end
				if(in == 4) begin
					state<=2268;
					out<=53;
				end
			end
			4158: begin
				if(in == 0) begin
					state<=4169;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=271;
					out<=56;
				end
				if(in == 3) begin
					state<=6158;
					out<=57;
				end
				if(in == 4) begin
					state<=2269;
					out<=58;
				end
			end
			4159: begin
				if(in == 0) begin
					state<=4170;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=272;
					out<=61;
				end
				if(in == 3) begin
					state<=6159;
					out<=62;
				end
				if(in == 4) begin
					state<=2270;
					out<=63;
				end
			end
			4160: begin
				if(in == 0) begin
					state<=4171;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=273;
					out<=66;
				end
				if(in == 3) begin
					state<=6160;
					out<=67;
				end
				if(in == 4) begin
					state<=2271;
					out<=68;
				end
			end
			4161: begin
				if(in == 0) begin
					state<=4172;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=274;
					out<=71;
				end
				if(in == 3) begin
					state<=6161;
					out<=72;
				end
				if(in == 4) begin
					state<=2272;
					out<=73;
				end
			end
			4162: begin
				if(in == 0) begin
					state<=4173;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=275;
					out<=76;
				end
				if(in == 3) begin
					state<=6162;
					out<=77;
				end
				if(in == 4) begin
					state<=2273;
					out<=78;
				end
			end
			4163: begin
				if(in == 0) begin
					state<=4174;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=276;
					out<=81;
				end
				if(in == 3) begin
					state<=6163;
					out<=82;
				end
				if(in == 4) begin
					state<=2274;
					out<=83;
				end
			end
			4164: begin
				if(in == 0) begin
					state<=4165;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=267;
					out<=86;
				end
				if(in == 3) begin
					state<=6154;
					out<=87;
				end
				if(in == 4) begin
					state<=2265;
					out<=88;
				end
			end
			4165: begin
				if(in == 0) begin
					state<=4176;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=278;
					out<=91;
				end
				if(in == 3) begin
					state<=6165;
					out<=92;
				end
				if(in == 4) begin
					state<=2276;
					out<=93;
				end
			end
			4166: begin
				if(in == 0) begin
					state<=4177;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=279;
					out<=96;
				end
				if(in == 3) begin
					state<=6166;
					out<=97;
				end
				if(in == 4) begin
					state<=2277;
					out<=98;
				end
			end
			4167: begin
				if(in == 0) begin
					state<=4178;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=280;
					out<=101;
				end
				if(in == 3) begin
					state<=6167;
					out<=102;
				end
				if(in == 4) begin
					state<=2278;
					out<=103;
				end
			end
			4168: begin
				if(in == 0) begin
					state<=4179;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=281;
					out<=106;
				end
				if(in == 3) begin
					state<=6168;
					out<=107;
				end
				if(in == 4) begin
					state<=2279;
					out<=108;
				end
			end
			4169: begin
				if(in == 0) begin
					state<=4180;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=282;
					out<=111;
				end
				if(in == 3) begin
					state<=6169;
					out<=112;
				end
				if(in == 4) begin
					state<=2280;
					out<=113;
				end
			end
			4170: begin
				if(in == 0) begin
					state<=4181;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=283;
					out<=116;
				end
				if(in == 3) begin
					state<=6170;
					out<=117;
				end
				if(in == 4) begin
					state<=2281;
					out<=118;
				end
			end
			4171: begin
				if(in == 0) begin
					state<=4182;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=284;
					out<=121;
				end
				if(in == 3) begin
					state<=6171;
					out<=122;
				end
				if(in == 4) begin
					state<=2282;
					out<=123;
				end
			end
			4172: begin
				if(in == 0) begin
					state<=4183;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=285;
					out<=126;
				end
				if(in == 3) begin
					state<=6172;
					out<=127;
				end
				if(in == 4) begin
					state<=2283;
					out<=128;
				end
			end
			4173: begin
				if(in == 0) begin
					state<=4184;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=286;
					out<=131;
				end
				if(in == 3) begin
					state<=6173;
					out<=132;
				end
				if(in == 4) begin
					state<=2284;
					out<=133;
				end
			end
			4174: begin
				if(in == 0) begin
					state<=4175;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=277;
					out<=136;
				end
				if(in == 3) begin
					state<=6164;
					out<=137;
				end
				if(in == 4) begin
					state<=2275;
					out<=138;
				end
			end
			4175: begin
				if(in == 0) begin
					state<=4186;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=288;
					out<=141;
				end
				if(in == 3) begin
					state<=6175;
					out<=142;
				end
				if(in == 4) begin
					state<=2286;
					out<=143;
				end
			end
			4176: begin
				if(in == 0) begin
					state<=4187;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=289;
					out<=146;
				end
				if(in == 3) begin
					state<=6176;
					out<=147;
				end
				if(in == 4) begin
					state<=2287;
					out<=148;
				end
			end
			4177: begin
				if(in == 0) begin
					state<=4188;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=290;
					out<=151;
				end
				if(in == 3) begin
					state<=6177;
					out<=152;
				end
				if(in == 4) begin
					state<=2288;
					out<=153;
				end
			end
			4178: begin
				if(in == 0) begin
					state<=4189;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=291;
					out<=156;
				end
				if(in == 3) begin
					state<=6178;
					out<=157;
				end
				if(in == 4) begin
					state<=2289;
					out<=158;
				end
			end
			4179: begin
				if(in == 0) begin
					state<=4190;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=292;
					out<=161;
				end
				if(in == 3) begin
					state<=6179;
					out<=162;
				end
				if(in == 4) begin
					state<=2290;
					out<=163;
				end
			end
			4180: begin
				if(in == 0) begin
					state<=4191;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=293;
					out<=166;
				end
				if(in == 3) begin
					state<=6180;
					out<=167;
				end
				if(in == 4) begin
					state<=2291;
					out<=168;
				end
			end
			4181: begin
				if(in == 0) begin
					state<=4192;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=294;
					out<=171;
				end
				if(in == 3) begin
					state<=6181;
					out<=172;
				end
				if(in == 4) begin
					state<=2292;
					out<=173;
				end
			end
			4182: begin
				if(in == 0) begin
					state<=4193;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=295;
					out<=176;
				end
				if(in == 3) begin
					state<=6182;
					out<=177;
				end
				if(in == 4) begin
					state<=2293;
					out<=178;
				end
			end
			4183: begin
				if(in == 0) begin
					state<=4194;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=296;
					out<=181;
				end
				if(in == 3) begin
					state<=6183;
					out<=182;
				end
				if(in == 4) begin
					state<=2294;
					out<=183;
				end
			end
			4184: begin
				if(in == 0) begin
					state<=4185;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=287;
					out<=186;
				end
				if(in == 3) begin
					state<=6174;
					out<=187;
				end
				if(in == 4) begin
					state<=2285;
					out<=188;
				end
			end
			4185: begin
				if(in == 0) begin
					state<=4196;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=298;
					out<=191;
				end
				if(in == 3) begin
					state<=6185;
					out<=192;
				end
				if(in == 4) begin
					state<=2296;
					out<=193;
				end
			end
			4186: begin
				if(in == 0) begin
					state<=4197;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=299;
					out<=196;
				end
				if(in == 3) begin
					state<=6186;
					out<=197;
				end
				if(in == 4) begin
					state<=2297;
					out<=198;
				end
			end
			4187: begin
				if(in == 0) begin
					state<=4198;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=300;
					out<=201;
				end
				if(in == 3) begin
					state<=6187;
					out<=202;
				end
				if(in == 4) begin
					state<=2298;
					out<=203;
				end
			end
			4188: begin
				if(in == 0) begin
					state<=4199;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=301;
					out<=206;
				end
				if(in == 3) begin
					state<=6188;
					out<=207;
				end
				if(in == 4) begin
					state<=2299;
					out<=208;
				end
			end
			4189: begin
				if(in == 0) begin
					state<=4200;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=302;
					out<=211;
				end
				if(in == 3) begin
					state<=6189;
					out<=212;
				end
				if(in == 4) begin
					state<=2300;
					out<=213;
				end
			end
			4190: begin
				if(in == 0) begin
					state<=4201;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=303;
					out<=216;
				end
				if(in == 3) begin
					state<=6190;
					out<=217;
				end
				if(in == 4) begin
					state<=2301;
					out<=218;
				end
			end
			4191: begin
				if(in == 0) begin
					state<=4202;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=304;
					out<=221;
				end
				if(in == 3) begin
					state<=6191;
					out<=222;
				end
				if(in == 4) begin
					state<=2302;
					out<=223;
				end
			end
			4192: begin
				if(in == 0) begin
					state<=4203;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=305;
					out<=226;
				end
				if(in == 3) begin
					state<=6192;
					out<=227;
				end
				if(in == 4) begin
					state<=2303;
					out<=228;
				end
			end
			4193: begin
				if(in == 0) begin
					state<=4204;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=306;
					out<=231;
				end
				if(in == 3) begin
					state<=6193;
					out<=232;
				end
				if(in == 4) begin
					state<=2304;
					out<=233;
				end
			end
			4194: begin
				if(in == 0) begin
					state<=4195;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=297;
					out<=236;
				end
				if(in == 3) begin
					state<=6184;
					out<=237;
				end
				if(in == 4) begin
					state<=2295;
					out<=238;
				end
			end
			4195: begin
				if(in == 0) begin
					state<=4206;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=308;
					out<=241;
				end
				if(in == 3) begin
					state<=6195;
					out<=242;
				end
				if(in == 4) begin
					state<=2306;
					out<=243;
				end
			end
			4196: begin
				if(in == 0) begin
					state<=4207;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=309;
					out<=246;
				end
				if(in == 3) begin
					state<=6196;
					out<=247;
				end
				if(in == 4) begin
					state<=2307;
					out<=248;
				end
			end
			4197: begin
				if(in == 0) begin
					state<=4208;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=310;
					out<=251;
				end
				if(in == 3) begin
					state<=6197;
					out<=252;
				end
				if(in == 4) begin
					state<=2308;
					out<=253;
				end
			end
			4198: begin
				if(in == 0) begin
					state<=4209;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=311;
					out<=0;
				end
				if(in == 3) begin
					state<=6198;
					out<=1;
				end
				if(in == 4) begin
					state<=2309;
					out<=2;
				end
			end
			4199: begin
				if(in == 0) begin
					state<=4210;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=312;
					out<=5;
				end
				if(in == 3) begin
					state<=6199;
					out<=6;
				end
				if(in == 4) begin
					state<=2310;
					out<=7;
				end
			end
			4200: begin
				if(in == 0) begin
					state<=4211;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=313;
					out<=10;
				end
				if(in == 3) begin
					state<=6200;
					out<=11;
				end
				if(in == 4) begin
					state<=2311;
					out<=12;
				end
			end
			4201: begin
				if(in == 0) begin
					state<=4212;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=314;
					out<=15;
				end
				if(in == 3) begin
					state<=6201;
					out<=16;
				end
				if(in == 4) begin
					state<=2312;
					out<=17;
				end
			end
			4202: begin
				if(in == 0) begin
					state<=4213;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=315;
					out<=20;
				end
				if(in == 3) begin
					state<=6202;
					out<=21;
				end
				if(in == 4) begin
					state<=2313;
					out<=22;
				end
			end
			4203: begin
				if(in == 0) begin
					state<=4214;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=316;
					out<=25;
				end
				if(in == 3) begin
					state<=6203;
					out<=26;
				end
				if(in == 4) begin
					state<=2314;
					out<=27;
				end
			end
			4204: begin
				if(in == 0) begin
					state<=4205;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=307;
					out<=30;
				end
				if(in == 3) begin
					state<=6194;
					out<=31;
				end
				if(in == 4) begin
					state<=2305;
					out<=32;
				end
			end
			4205: begin
				if(in == 0) begin
					state<=4216;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=318;
					out<=35;
				end
				if(in == 3) begin
					state<=6205;
					out<=36;
				end
				if(in == 4) begin
					state<=2316;
					out<=37;
				end
			end
			4206: begin
				if(in == 0) begin
					state<=4217;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=319;
					out<=40;
				end
				if(in == 3) begin
					state<=6206;
					out<=41;
				end
				if(in == 4) begin
					state<=2317;
					out<=42;
				end
			end
			4207: begin
				if(in == 0) begin
					state<=4218;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=320;
					out<=45;
				end
				if(in == 3) begin
					state<=6207;
					out<=46;
				end
				if(in == 4) begin
					state<=2318;
					out<=47;
				end
			end
			4208: begin
				if(in == 0) begin
					state<=4219;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=321;
					out<=50;
				end
				if(in == 3) begin
					state<=6208;
					out<=51;
				end
				if(in == 4) begin
					state<=2319;
					out<=52;
				end
			end
			4209: begin
				if(in == 0) begin
					state<=4220;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=322;
					out<=55;
				end
				if(in == 3) begin
					state<=6209;
					out<=56;
				end
				if(in == 4) begin
					state<=2320;
					out<=57;
				end
			end
			4210: begin
				if(in == 0) begin
					state<=4221;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=323;
					out<=60;
				end
				if(in == 3) begin
					state<=6210;
					out<=61;
				end
				if(in == 4) begin
					state<=2321;
					out<=62;
				end
			end
			4211: begin
				if(in == 0) begin
					state<=4222;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=324;
					out<=65;
				end
				if(in == 3) begin
					state<=6211;
					out<=66;
				end
				if(in == 4) begin
					state<=2322;
					out<=67;
				end
			end
			4212: begin
				if(in == 0) begin
					state<=4223;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=325;
					out<=70;
				end
				if(in == 3) begin
					state<=6212;
					out<=71;
				end
				if(in == 4) begin
					state<=2323;
					out<=72;
				end
			end
			4213: begin
				if(in == 0) begin
					state<=4224;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=326;
					out<=75;
				end
				if(in == 3) begin
					state<=6213;
					out<=76;
				end
				if(in == 4) begin
					state<=2324;
					out<=77;
				end
			end
			4214: begin
				if(in == 0) begin
					state<=4215;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=317;
					out<=80;
				end
				if(in == 3) begin
					state<=6204;
					out<=81;
				end
				if(in == 4) begin
					state<=2315;
					out<=82;
				end
			end
			4215: begin
				if(in == 0) begin
					state<=5343;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=1454;
					out<=85;
				end
				if(in == 3) begin
					state<=6788;
					out<=86;
				end
				if(in == 4) begin
					state<=2899;
					out<=87;
				end
			end
			4216: begin
				if(in == 0) begin
					state<=5344;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=1455;
					out<=90;
				end
				if(in == 3) begin
					state<=6789;
					out<=91;
				end
				if(in == 4) begin
					state<=2900;
					out<=92;
				end
			end
			4217: begin
				if(in == 0) begin
					state<=5345;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=1456;
					out<=95;
				end
				if(in == 3) begin
					state<=6790;
					out<=96;
				end
				if(in == 4) begin
					state<=2901;
					out<=97;
				end
			end
			4218: begin
				if(in == 0) begin
					state<=5346;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=1457;
					out<=100;
				end
				if(in == 3) begin
					state<=6791;
					out<=101;
				end
				if(in == 4) begin
					state<=2902;
					out<=102;
				end
			end
			4219: begin
				if(in == 0) begin
					state<=5347;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=1458;
					out<=105;
				end
				if(in == 3) begin
					state<=6792;
					out<=106;
				end
				if(in == 4) begin
					state<=2903;
					out<=107;
				end
			end
			4220: begin
				if(in == 0) begin
					state<=5348;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=1459;
					out<=110;
				end
				if(in == 3) begin
					state<=6793;
					out<=111;
				end
				if(in == 4) begin
					state<=2904;
					out<=112;
				end
			end
			4221: begin
				if(in == 0) begin
					state<=5349;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=1460;
					out<=115;
				end
				if(in == 3) begin
					state<=6794;
					out<=116;
				end
				if(in == 4) begin
					state<=2905;
					out<=117;
				end
			end
			4222: begin
				if(in == 0) begin
					state<=5350;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=1461;
					out<=120;
				end
				if(in == 3) begin
					state<=6795;
					out<=121;
				end
				if(in == 4) begin
					state<=2906;
					out<=122;
				end
			end
			4223: begin
				if(in == 0) begin
					state<=5351;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=1462;
					out<=125;
				end
				if(in == 3) begin
					state<=6796;
					out<=126;
				end
				if(in == 4) begin
					state<=2907;
					out<=127;
				end
			end
			4224: begin
				if(in == 0) begin
					state<=5342;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=1453;
					out<=130;
				end
				if(in == 3) begin
					state<=6787;
					out<=131;
				end
				if(in == 4) begin
					state<=2898;
					out<=132;
				end
			end
			4225: begin
				if(in == 0) begin
					state<=4236;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=338;
					out<=135;
				end
				if(in == 3) begin
					state<=6225;
					out<=136;
				end
				if(in == 4) begin
					state<=2336;
					out<=137;
				end
			end
			4226: begin
				if(in == 0) begin
					state<=4237;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=339;
					out<=140;
				end
				if(in == 3) begin
					state<=6226;
					out<=141;
				end
				if(in == 4) begin
					state<=2337;
					out<=142;
				end
			end
			4227: begin
				if(in == 0) begin
					state<=4238;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=340;
					out<=145;
				end
				if(in == 3) begin
					state<=6227;
					out<=146;
				end
				if(in == 4) begin
					state<=2338;
					out<=147;
				end
			end
			4228: begin
				if(in == 0) begin
					state<=4239;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=341;
					out<=150;
				end
				if(in == 3) begin
					state<=6228;
					out<=151;
				end
				if(in == 4) begin
					state<=2339;
					out<=152;
				end
			end
			4229: begin
				if(in == 0) begin
					state<=4240;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=342;
					out<=155;
				end
				if(in == 3) begin
					state<=6229;
					out<=156;
				end
				if(in == 4) begin
					state<=2340;
					out<=157;
				end
			end
			4230: begin
				if(in == 0) begin
					state<=4241;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=343;
					out<=160;
				end
				if(in == 3) begin
					state<=6230;
					out<=161;
				end
				if(in == 4) begin
					state<=2341;
					out<=162;
				end
			end
			4231: begin
				if(in == 0) begin
					state<=4242;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=344;
					out<=165;
				end
				if(in == 3) begin
					state<=6231;
					out<=166;
				end
				if(in == 4) begin
					state<=2342;
					out<=167;
				end
			end
			4232: begin
				if(in == 0) begin
					state<=4243;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=345;
					out<=170;
				end
				if(in == 3) begin
					state<=6232;
					out<=171;
				end
				if(in == 4) begin
					state<=2343;
					out<=172;
				end
			end
			4233: begin
				if(in == 0) begin
					state<=4234;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=336;
					out<=175;
				end
				if(in == 3) begin
					state<=6223;
					out<=176;
				end
				if(in == 4) begin
					state<=2334;
					out<=177;
				end
			end
			4234: begin
				if(in == 0) begin
					state<=4245;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=347;
					out<=180;
				end
				if(in == 3) begin
					state<=6234;
					out<=181;
				end
				if(in == 4) begin
					state<=2345;
					out<=182;
				end
			end
			4235: begin
				if(in == 0) begin
					state<=4246;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=348;
					out<=185;
				end
				if(in == 3) begin
					state<=6235;
					out<=186;
				end
				if(in == 4) begin
					state<=2346;
					out<=187;
				end
			end
			4236: begin
				if(in == 0) begin
					state<=4247;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=349;
					out<=190;
				end
				if(in == 3) begin
					state<=6236;
					out<=191;
				end
				if(in == 4) begin
					state<=2347;
					out<=192;
				end
			end
			4237: begin
				if(in == 0) begin
					state<=4248;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=350;
					out<=195;
				end
				if(in == 3) begin
					state<=6237;
					out<=196;
				end
				if(in == 4) begin
					state<=2348;
					out<=197;
				end
			end
			4238: begin
				if(in == 0) begin
					state<=4249;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=351;
					out<=200;
				end
				if(in == 3) begin
					state<=6238;
					out<=201;
				end
				if(in == 4) begin
					state<=2349;
					out<=202;
				end
			end
			4239: begin
				if(in == 0) begin
					state<=4250;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=352;
					out<=205;
				end
				if(in == 3) begin
					state<=6239;
					out<=206;
				end
				if(in == 4) begin
					state<=2350;
					out<=207;
				end
			end
			4240: begin
				if(in == 0) begin
					state<=4251;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=353;
					out<=210;
				end
				if(in == 3) begin
					state<=6240;
					out<=211;
				end
				if(in == 4) begin
					state<=2351;
					out<=212;
				end
			end
			4241: begin
				if(in == 0) begin
					state<=4252;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=354;
					out<=215;
				end
				if(in == 3) begin
					state<=6241;
					out<=216;
				end
				if(in == 4) begin
					state<=2352;
					out<=217;
				end
			end
			4242: begin
				if(in == 0) begin
					state<=4253;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=355;
					out<=220;
				end
				if(in == 3) begin
					state<=6242;
					out<=221;
				end
				if(in == 4) begin
					state<=2353;
					out<=222;
				end
			end
			4243: begin
				if(in == 0) begin
					state<=4244;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=346;
					out<=225;
				end
				if(in == 3) begin
					state<=6233;
					out<=226;
				end
				if(in == 4) begin
					state<=2344;
					out<=227;
				end
			end
			4244: begin
				if(in == 0) begin
					state<=4255;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=357;
					out<=230;
				end
				if(in == 3) begin
					state<=6829;
					out<=231;
				end
				if(in == 4) begin
					state<=2940;
					out<=232;
				end
			end
			4245: begin
				if(in == 0) begin
					state<=4256;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=358;
					out<=235;
				end
				if(in == 3) begin
					state<=6830;
					out<=236;
				end
				if(in == 4) begin
					state<=2941;
					out<=237;
				end
			end
			4246: begin
				if(in == 0) begin
					state<=4257;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=359;
					out<=240;
				end
				if(in == 3) begin
					state<=6831;
					out<=241;
				end
				if(in == 4) begin
					state<=2942;
					out<=242;
				end
			end
			4247: begin
				if(in == 0) begin
					state<=4258;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=360;
					out<=245;
				end
				if(in == 3) begin
					state<=6832;
					out<=246;
				end
				if(in == 4) begin
					state<=2943;
					out<=247;
				end
			end
			4248: begin
				if(in == 0) begin
					state<=4259;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=361;
					out<=250;
				end
				if(in == 3) begin
					state<=6833;
					out<=251;
				end
				if(in == 4) begin
					state<=2944;
					out<=252;
				end
			end
			4249: begin
				if(in == 0) begin
					state<=4260;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=362;
					out<=255;
				end
				if(in == 3) begin
					state<=6834;
					out<=0;
				end
				if(in == 4) begin
					state<=2945;
					out<=1;
				end
			end
			4250: begin
				if(in == 0) begin
					state<=4261;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=363;
					out<=4;
				end
				if(in == 3) begin
					state<=6835;
					out<=5;
				end
				if(in == 4) begin
					state<=2946;
					out<=6;
				end
			end
			4251: begin
				if(in == 0) begin
					state<=4262;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=364;
					out<=9;
				end
				if(in == 3) begin
					state<=6836;
					out<=10;
				end
				if(in == 4) begin
					state<=2947;
					out<=11;
				end
			end
			4252: begin
				if(in == 0) begin
					state<=4263;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=365;
					out<=14;
				end
				if(in == 3) begin
					state<=6837;
					out<=15;
				end
				if(in == 4) begin
					state<=2948;
					out<=16;
				end
			end
			4253: begin
				if(in == 0) begin
					state<=4254;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=356;
					out<=19;
				end
				if(in == 3) begin
					state<=6828;
					out<=20;
				end
				if(in == 4) begin
					state<=2939;
					out<=21;
				end
			end
			4254: begin
				if(in == 0) begin
					state<=4265;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=367;
					out<=24;
				end
				if(in == 3) begin
					state<=6839;
					out<=25;
				end
				if(in == 4) begin
					state<=2950;
					out<=26;
				end
			end
			4255: begin
				if(in == 0) begin
					state<=4266;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=368;
					out<=29;
				end
				if(in == 3) begin
					state<=6840;
					out<=30;
				end
				if(in == 4) begin
					state<=2951;
					out<=31;
				end
			end
			4256: begin
				if(in == 0) begin
					state<=4267;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=369;
					out<=34;
				end
				if(in == 3) begin
					state<=6841;
					out<=35;
				end
				if(in == 4) begin
					state<=2952;
					out<=36;
				end
			end
			4257: begin
				if(in == 0) begin
					state<=4268;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=370;
					out<=39;
				end
				if(in == 3) begin
					state<=6842;
					out<=40;
				end
				if(in == 4) begin
					state<=2953;
					out<=41;
				end
			end
			4258: begin
				if(in == 0) begin
					state<=4269;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=371;
					out<=44;
				end
				if(in == 3) begin
					state<=6843;
					out<=45;
				end
				if(in == 4) begin
					state<=2954;
					out<=46;
				end
			end
			4259: begin
				if(in == 0) begin
					state<=4270;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=372;
					out<=49;
				end
				if(in == 3) begin
					state<=6844;
					out<=50;
				end
				if(in == 4) begin
					state<=2955;
					out<=51;
				end
			end
			4260: begin
				if(in == 0) begin
					state<=4271;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=373;
					out<=54;
				end
				if(in == 3) begin
					state<=6845;
					out<=55;
				end
				if(in == 4) begin
					state<=2956;
					out<=56;
				end
			end
			4261: begin
				if(in == 0) begin
					state<=4272;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=374;
					out<=59;
				end
				if(in == 3) begin
					state<=6846;
					out<=60;
				end
				if(in == 4) begin
					state<=2957;
					out<=61;
				end
			end
			4262: begin
				if(in == 0) begin
					state<=4273;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=375;
					out<=64;
				end
				if(in == 3) begin
					state<=6847;
					out<=65;
				end
				if(in == 4) begin
					state<=2958;
					out<=66;
				end
			end
			4263: begin
				if(in == 0) begin
					state<=4264;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=366;
					out<=69;
				end
				if(in == 3) begin
					state<=6838;
					out<=70;
				end
				if(in == 4) begin
					state<=2949;
					out<=71;
				end
			end
			4264: begin
				if(in == 0) begin
					state<=4275;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=377;
					out<=74;
				end
				if(in == 3) begin
					state<=6849;
					out<=75;
				end
				if(in == 4) begin
					state<=2960;
					out<=76;
				end
			end
			4265: begin
				if(in == 0) begin
					state<=4276;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=378;
					out<=79;
				end
				if(in == 3) begin
					state<=6850;
					out<=80;
				end
				if(in == 4) begin
					state<=2961;
					out<=81;
				end
			end
			4266: begin
				if(in == 0) begin
					state<=4277;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=379;
					out<=84;
				end
				if(in == 3) begin
					state<=6851;
					out<=85;
				end
				if(in == 4) begin
					state<=2962;
					out<=86;
				end
			end
			4267: begin
				if(in == 0) begin
					state<=4278;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=380;
					out<=89;
				end
				if(in == 3) begin
					state<=6852;
					out<=90;
				end
				if(in == 4) begin
					state<=2963;
					out<=91;
				end
			end
			4268: begin
				if(in == 0) begin
					state<=4279;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=381;
					out<=94;
				end
				if(in == 3) begin
					state<=6853;
					out<=95;
				end
				if(in == 4) begin
					state<=2964;
					out<=96;
				end
			end
			4269: begin
				if(in == 0) begin
					state<=4280;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=382;
					out<=99;
				end
				if(in == 3) begin
					state<=6854;
					out<=100;
				end
				if(in == 4) begin
					state<=2965;
					out<=101;
				end
			end
			4270: begin
				if(in == 0) begin
					state<=4281;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=383;
					out<=104;
				end
				if(in == 3) begin
					state<=6855;
					out<=105;
				end
				if(in == 4) begin
					state<=2966;
					out<=106;
				end
			end
			4271: begin
				if(in == 0) begin
					state<=4282;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=384;
					out<=109;
				end
				if(in == 3) begin
					state<=6856;
					out<=110;
				end
				if(in == 4) begin
					state<=2967;
					out<=111;
				end
			end
			4272: begin
				if(in == 0) begin
					state<=4283;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=385;
					out<=114;
				end
				if(in == 3) begin
					state<=6857;
					out<=115;
				end
				if(in == 4) begin
					state<=2968;
					out<=116;
				end
			end
			4273: begin
				if(in == 0) begin
					state<=4274;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=376;
					out<=119;
				end
				if(in == 3) begin
					state<=6848;
					out<=120;
				end
				if(in == 4) begin
					state<=2959;
					out<=121;
				end
			end
			4274: begin
				if(in == 0) begin
					state<=4285;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=387;
					out<=124;
				end
				if(in == 3) begin
					state<=6859;
					out<=125;
				end
				if(in == 4) begin
					state<=2970;
					out<=126;
				end
			end
			4275: begin
				if(in == 0) begin
					state<=4286;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=388;
					out<=129;
				end
				if(in == 3) begin
					state<=6860;
					out<=130;
				end
				if(in == 4) begin
					state<=2971;
					out<=131;
				end
			end
			4276: begin
				if(in == 0) begin
					state<=4287;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=389;
					out<=134;
				end
				if(in == 3) begin
					state<=6861;
					out<=135;
				end
				if(in == 4) begin
					state<=2972;
					out<=136;
				end
			end
			4277: begin
				if(in == 0) begin
					state<=4288;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=390;
					out<=139;
				end
				if(in == 3) begin
					state<=6862;
					out<=140;
				end
				if(in == 4) begin
					state<=2973;
					out<=141;
				end
			end
			4278: begin
				if(in == 0) begin
					state<=4289;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=391;
					out<=144;
				end
				if(in == 3) begin
					state<=6863;
					out<=145;
				end
				if(in == 4) begin
					state<=2974;
					out<=146;
				end
			end
			4279: begin
				if(in == 0) begin
					state<=4290;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=392;
					out<=149;
				end
				if(in == 3) begin
					state<=6864;
					out<=150;
				end
				if(in == 4) begin
					state<=2975;
					out<=151;
				end
			end
			4280: begin
				if(in == 0) begin
					state<=4291;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=393;
					out<=154;
				end
				if(in == 3) begin
					state<=6865;
					out<=155;
				end
				if(in == 4) begin
					state<=2976;
					out<=156;
				end
			end
			4281: begin
				if(in == 0) begin
					state<=4292;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=394;
					out<=159;
				end
				if(in == 3) begin
					state<=6866;
					out<=160;
				end
				if(in == 4) begin
					state<=2977;
					out<=161;
				end
			end
			4282: begin
				if(in == 0) begin
					state<=4293;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=395;
					out<=164;
				end
				if(in == 3) begin
					state<=6867;
					out<=165;
				end
				if(in == 4) begin
					state<=2978;
					out<=166;
				end
			end
			4283: begin
				if(in == 0) begin
					state<=4284;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=386;
					out<=169;
				end
				if(in == 3) begin
					state<=6858;
					out<=170;
				end
				if(in == 4) begin
					state<=2969;
					out<=171;
				end
			end
			4284: begin
				if(in == 0) begin
					state<=4898;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=1000;
					out<=174;
				end
				if(in == 3) begin
					state<=6869;
					out<=175;
				end
				if(in == 4) begin
					state<=2980;
					out<=176;
				end
			end
			4285: begin
				if(in == 0) begin
					state<=4899;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=1001;
					out<=179;
				end
				if(in == 3) begin
					state<=6870;
					out<=180;
				end
				if(in == 4) begin
					state<=2981;
					out<=181;
				end
			end
			4286: begin
				if(in == 0) begin
					state<=4900;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=1002;
					out<=184;
				end
				if(in == 3) begin
					state<=6871;
					out<=185;
				end
				if(in == 4) begin
					state<=2982;
					out<=186;
				end
			end
			4287: begin
				if(in == 0) begin
					state<=4901;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=1003;
					out<=189;
				end
				if(in == 3) begin
					state<=6872;
					out<=190;
				end
				if(in == 4) begin
					state<=2983;
					out<=191;
				end
			end
			4288: begin
				if(in == 0) begin
					state<=4902;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=1004;
					out<=194;
				end
				if(in == 3) begin
					state<=6873;
					out<=195;
				end
				if(in == 4) begin
					state<=2984;
					out<=196;
				end
			end
			4289: begin
				if(in == 0) begin
					state<=4903;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=1005;
					out<=199;
				end
				if(in == 3) begin
					state<=6874;
					out<=200;
				end
				if(in == 4) begin
					state<=2985;
					out<=201;
				end
			end
			4290: begin
				if(in == 0) begin
					state<=4904;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=1006;
					out<=204;
				end
				if(in == 3) begin
					state<=6875;
					out<=205;
				end
				if(in == 4) begin
					state<=2986;
					out<=206;
				end
			end
			4291: begin
				if(in == 0) begin
					state<=4905;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=1007;
					out<=209;
				end
				if(in == 3) begin
					state<=6876;
					out<=210;
				end
				if(in == 4) begin
					state<=2987;
					out<=211;
				end
			end
			4292: begin
				if(in == 0) begin
					state<=4906;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=1008;
					out<=214;
				end
				if(in == 3) begin
					state<=6877;
					out<=215;
				end
				if(in == 4) begin
					state<=2988;
					out<=216;
				end
			end
			4293: begin
				if(in == 0) begin
					state<=4897;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=999;
					out<=219;
				end
				if(in == 3) begin
					state<=6868;
					out<=220;
				end
				if(in == 4) begin
					state<=2979;
					out<=221;
				end
			end
			4294: begin
				if(in == 0) begin
					state<=4305;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=407;
					out<=224;
				end
				if(in == 3) begin
					state<=6910;
					out<=225;
				end
				if(in == 4) begin
					state<=3021;
					out<=226;
				end
			end
			4295: begin
				if(in == 0) begin
					state<=4306;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=408;
					out<=229;
				end
				if(in == 3) begin
					state<=6911;
					out<=230;
				end
				if(in == 4) begin
					state<=3022;
					out<=231;
				end
			end
			4296: begin
				if(in == 0) begin
					state<=4307;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=409;
					out<=234;
				end
				if(in == 3) begin
					state<=6912;
					out<=235;
				end
				if(in == 4) begin
					state<=3023;
					out<=236;
				end
			end
			4297: begin
				if(in == 0) begin
					state<=4308;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=410;
					out<=239;
				end
				if(in == 3) begin
					state<=6913;
					out<=240;
				end
				if(in == 4) begin
					state<=3024;
					out<=241;
				end
			end
			4298: begin
				if(in == 0) begin
					state<=4309;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=411;
					out<=244;
				end
				if(in == 3) begin
					state<=6914;
					out<=245;
				end
				if(in == 4) begin
					state<=3025;
					out<=246;
				end
			end
			4299: begin
				if(in == 0) begin
					state<=4310;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=412;
					out<=249;
				end
				if(in == 3) begin
					state<=6915;
					out<=250;
				end
				if(in == 4) begin
					state<=3026;
					out<=251;
				end
			end
			4300: begin
				if(in == 0) begin
					state<=4311;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=413;
					out<=254;
				end
				if(in == 3) begin
					state<=6916;
					out<=255;
				end
				if(in == 4) begin
					state<=3027;
					out<=0;
				end
			end
			4301: begin
				if(in == 0) begin
					state<=4312;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=414;
					out<=3;
				end
				if(in == 3) begin
					state<=6917;
					out<=4;
				end
				if(in == 4) begin
					state<=3028;
					out<=5;
				end
			end
			4302: begin
				if(in == 0) begin
					state<=4303;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=405;
					out<=8;
				end
				if(in == 3) begin
					state<=6908;
					out<=9;
				end
				if(in == 4) begin
					state<=3019;
					out<=10;
				end
			end
			4303: begin
				if(in == 0) begin
					state<=4929;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=1031;
					out<=13;
				end
				if(in == 3) begin
					state<=6919;
					out<=14;
				end
				if(in == 4) begin
					state<=3030;
					out<=15;
				end
			end
			4304: begin
				if(in == 0) begin
					state<=4930;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=1032;
					out<=18;
				end
				if(in == 3) begin
					state<=6920;
					out<=19;
				end
				if(in == 4) begin
					state<=3031;
					out<=20;
				end
			end
			4305: begin
				if(in == 0) begin
					state<=4931;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=1033;
					out<=23;
				end
				if(in == 3) begin
					state<=6921;
					out<=24;
				end
				if(in == 4) begin
					state<=3032;
					out<=25;
				end
			end
			4306: begin
				if(in == 0) begin
					state<=4932;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=1034;
					out<=28;
				end
				if(in == 3) begin
					state<=6922;
					out<=29;
				end
				if(in == 4) begin
					state<=3033;
					out<=30;
				end
			end
			4307: begin
				if(in == 0) begin
					state<=4933;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=1035;
					out<=33;
				end
				if(in == 3) begin
					state<=6923;
					out<=34;
				end
				if(in == 4) begin
					state<=3034;
					out<=35;
				end
			end
			4308: begin
				if(in == 0) begin
					state<=4934;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=1036;
					out<=38;
				end
				if(in == 3) begin
					state<=6924;
					out<=39;
				end
				if(in == 4) begin
					state<=3035;
					out<=40;
				end
			end
			4309: begin
				if(in == 0) begin
					state<=4935;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=1037;
					out<=43;
				end
				if(in == 3) begin
					state<=6925;
					out<=44;
				end
				if(in == 4) begin
					state<=3036;
					out<=45;
				end
			end
			4310: begin
				if(in == 0) begin
					state<=4936;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=1038;
					out<=48;
				end
				if(in == 3) begin
					state<=6926;
					out<=49;
				end
				if(in == 4) begin
					state<=3037;
					out<=50;
				end
			end
			4311: begin
				if(in == 0) begin
					state<=4937;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=1039;
					out<=53;
				end
				if(in == 3) begin
					state<=6927;
					out<=54;
				end
				if(in == 4) begin
					state<=3038;
					out<=55;
				end
			end
			4312: begin
				if(in == 0) begin
					state<=4928;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=1030;
					out<=58;
				end
				if(in == 3) begin
					state<=6918;
					out<=59;
				end
				if(in == 4) begin
					state<=3029;
					out<=60;
				end
			end
			4313: begin
				if(in == 0) begin
					state<=4324;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=426;
					out<=63;
				end
				if(in == 3) begin
					state<=6313;
					out<=64;
				end
				if(in == 4) begin
					state<=2424;
					out<=65;
				end
			end
			4314: begin
				if(in == 0) begin
					state<=4325;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=427;
					out<=68;
				end
				if(in == 3) begin
					state<=6314;
					out<=69;
				end
				if(in == 4) begin
					state<=2425;
					out<=70;
				end
			end
			4315: begin
				if(in == 0) begin
					state<=4326;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=428;
					out<=73;
				end
				if(in == 3) begin
					state<=6315;
					out<=74;
				end
				if(in == 4) begin
					state<=2426;
					out<=75;
				end
			end
			4316: begin
				if(in == 0) begin
					state<=4327;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=429;
					out<=78;
				end
				if(in == 3) begin
					state<=6316;
					out<=79;
				end
				if(in == 4) begin
					state<=2427;
					out<=80;
				end
			end
			4317: begin
				if(in == 0) begin
					state<=4328;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=430;
					out<=83;
				end
				if(in == 3) begin
					state<=6317;
					out<=84;
				end
				if(in == 4) begin
					state<=2428;
					out<=85;
				end
			end
			4318: begin
				if(in == 0) begin
					state<=4329;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=431;
					out<=88;
				end
				if(in == 3) begin
					state<=6318;
					out<=89;
				end
				if(in == 4) begin
					state<=2429;
					out<=90;
				end
			end
			4319: begin
				if(in == 0) begin
					state<=4330;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=432;
					out<=93;
				end
				if(in == 3) begin
					state<=6319;
					out<=94;
				end
				if(in == 4) begin
					state<=2430;
					out<=95;
				end
			end
			4320: begin
				if(in == 0) begin
					state<=4331;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=433;
					out<=98;
				end
				if(in == 3) begin
					state<=6320;
					out<=99;
				end
				if(in == 4) begin
					state<=2431;
					out<=100;
				end
			end
			4321: begin
				if(in == 0) begin
					state<=4332;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=434;
					out<=103;
				end
				if(in == 3) begin
					state<=6321;
					out<=104;
				end
				if(in == 4) begin
					state<=2432;
					out<=105;
				end
			end
			4322: begin
				if(in == 0) begin
					state<=4323;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=425;
					out<=108;
				end
				if(in == 3) begin
					state<=6312;
					out<=109;
				end
				if(in == 4) begin
					state<=2423;
					out<=110;
				end
			end
			4323: begin
				if(in == 0) begin
					state<=4334;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=436;
					out<=113;
				end
				if(in == 3) begin
					state<=6323;
					out<=114;
				end
				if(in == 4) begin
					state<=2434;
					out<=115;
				end
			end
			4324: begin
				if(in == 0) begin
					state<=4335;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=437;
					out<=118;
				end
				if(in == 3) begin
					state<=6324;
					out<=119;
				end
				if(in == 4) begin
					state<=2435;
					out<=120;
				end
			end
			4325: begin
				if(in == 0) begin
					state<=4336;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=438;
					out<=123;
				end
				if(in == 3) begin
					state<=6325;
					out<=124;
				end
				if(in == 4) begin
					state<=2436;
					out<=125;
				end
			end
			4326: begin
				if(in == 0) begin
					state<=4337;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=439;
					out<=128;
				end
				if(in == 3) begin
					state<=6326;
					out<=129;
				end
				if(in == 4) begin
					state<=2437;
					out<=130;
				end
			end
			4327: begin
				if(in == 0) begin
					state<=4338;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=440;
					out<=133;
				end
				if(in == 3) begin
					state<=6327;
					out<=134;
				end
				if(in == 4) begin
					state<=2438;
					out<=135;
				end
			end
			4328: begin
				if(in == 0) begin
					state<=4339;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=441;
					out<=138;
				end
				if(in == 3) begin
					state<=6328;
					out<=139;
				end
				if(in == 4) begin
					state<=2439;
					out<=140;
				end
			end
			4329: begin
				if(in == 0) begin
					state<=4340;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=442;
					out<=143;
				end
				if(in == 3) begin
					state<=6329;
					out<=144;
				end
				if(in == 4) begin
					state<=2440;
					out<=145;
				end
			end
			4330: begin
				if(in == 0) begin
					state<=4341;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=443;
					out<=148;
				end
				if(in == 3) begin
					state<=6330;
					out<=149;
				end
				if(in == 4) begin
					state<=2441;
					out<=150;
				end
			end
			4331: begin
				if(in == 0) begin
					state<=4342;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=444;
					out<=153;
				end
				if(in == 3) begin
					state<=6331;
					out<=154;
				end
				if(in == 4) begin
					state<=2442;
					out<=155;
				end
			end
			4332: begin
				if(in == 0) begin
					state<=4333;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=435;
					out<=158;
				end
				if(in == 3) begin
					state<=6322;
					out<=159;
				end
				if(in == 4) begin
					state<=2433;
					out<=160;
				end
			end
			4333: begin
				if(in == 0) begin
					state<=4344;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=446;
					out<=163;
				end
				if(in == 3) begin
					state<=6333;
					out<=164;
				end
				if(in == 4) begin
					state<=2444;
					out<=165;
				end
			end
			4334: begin
				if(in == 0) begin
					state<=4345;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=447;
					out<=168;
				end
				if(in == 3) begin
					state<=6334;
					out<=169;
				end
				if(in == 4) begin
					state<=2445;
					out<=170;
				end
			end
			4335: begin
				if(in == 0) begin
					state<=4346;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=448;
					out<=173;
				end
				if(in == 3) begin
					state<=6335;
					out<=174;
				end
				if(in == 4) begin
					state<=2446;
					out<=175;
				end
			end
			4336: begin
				if(in == 0) begin
					state<=4347;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=449;
					out<=178;
				end
				if(in == 3) begin
					state<=6336;
					out<=179;
				end
				if(in == 4) begin
					state<=2447;
					out<=180;
				end
			end
			4337: begin
				if(in == 0) begin
					state<=4348;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=450;
					out<=183;
				end
				if(in == 3) begin
					state<=6337;
					out<=184;
				end
				if(in == 4) begin
					state<=2448;
					out<=185;
				end
			end
			4338: begin
				if(in == 0) begin
					state<=4349;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=451;
					out<=188;
				end
				if(in == 3) begin
					state<=6338;
					out<=189;
				end
				if(in == 4) begin
					state<=2449;
					out<=190;
				end
			end
			4339: begin
				if(in == 0) begin
					state<=4350;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=452;
					out<=193;
				end
				if(in == 3) begin
					state<=6339;
					out<=194;
				end
				if(in == 4) begin
					state<=2450;
					out<=195;
				end
			end
			4340: begin
				if(in == 0) begin
					state<=4351;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=453;
					out<=198;
				end
				if(in == 3) begin
					state<=6340;
					out<=199;
				end
				if(in == 4) begin
					state<=2451;
					out<=200;
				end
			end
			4341: begin
				if(in == 0) begin
					state<=4352;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=454;
					out<=203;
				end
				if(in == 3) begin
					state<=6341;
					out<=204;
				end
				if(in == 4) begin
					state<=2452;
					out<=205;
				end
			end
			4342: begin
				if(in == 0) begin
					state<=4343;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=445;
					out<=208;
				end
				if(in == 3) begin
					state<=6332;
					out<=209;
				end
				if(in == 4) begin
					state<=2443;
					out<=210;
				end
			end
			4343: begin
				if(in == 0) begin
					state<=4354;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=456;
					out<=213;
				end
				if(in == 3) begin
					state<=6343;
					out<=214;
				end
				if(in == 4) begin
					state<=2454;
					out<=215;
				end
			end
			4344: begin
				if(in == 0) begin
					state<=4355;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=457;
					out<=218;
				end
				if(in == 3) begin
					state<=6344;
					out<=219;
				end
				if(in == 4) begin
					state<=2455;
					out<=220;
				end
			end
			4345: begin
				if(in == 0) begin
					state<=4356;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=458;
					out<=223;
				end
				if(in == 3) begin
					state<=6345;
					out<=224;
				end
				if(in == 4) begin
					state<=2456;
					out<=225;
				end
			end
			4346: begin
				if(in == 0) begin
					state<=4357;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=459;
					out<=228;
				end
				if(in == 3) begin
					state<=6346;
					out<=229;
				end
				if(in == 4) begin
					state<=2457;
					out<=230;
				end
			end
			4347: begin
				if(in == 0) begin
					state<=4358;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=460;
					out<=233;
				end
				if(in == 3) begin
					state<=6347;
					out<=234;
				end
				if(in == 4) begin
					state<=2458;
					out<=235;
				end
			end
			4348: begin
				if(in == 0) begin
					state<=4359;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=461;
					out<=238;
				end
				if(in == 3) begin
					state<=6348;
					out<=239;
				end
				if(in == 4) begin
					state<=2459;
					out<=240;
				end
			end
			4349: begin
				if(in == 0) begin
					state<=4360;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=462;
					out<=243;
				end
				if(in == 3) begin
					state<=6349;
					out<=244;
				end
				if(in == 4) begin
					state<=2460;
					out<=245;
				end
			end
			4350: begin
				if(in == 0) begin
					state<=4361;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=463;
					out<=248;
				end
				if(in == 3) begin
					state<=6350;
					out<=249;
				end
				if(in == 4) begin
					state<=2461;
					out<=250;
				end
			end
			4351: begin
				if(in == 0) begin
					state<=4362;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=464;
					out<=253;
				end
				if(in == 3) begin
					state<=6351;
					out<=254;
				end
				if(in == 4) begin
					state<=2462;
					out<=255;
				end
			end
			4352: begin
				if(in == 0) begin
					state<=4353;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=455;
					out<=2;
				end
				if(in == 3) begin
					state<=6342;
					out<=3;
				end
				if(in == 4) begin
					state<=2453;
					out<=4;
				end
			end
			4353: begin
				if(in == 0) begin
					state<=5374;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=1485;
					out<=7;
				end
				if(in == 3) begin
					state<=7306;
					out<=8;
				end
				if(in == 4) begin
					state<=3417;
					out<=9;
				end
			end
			4354: begin
				if(in == 0) begin
					state<=5375;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=1486;
					out<=12;
				end
				if(in == 3) begin
					state<=7307;
					out<=13;
				end
				if(in == 4) begin
					state<=3418;
					out<=14;
				end
			end
			4355: begin
				if(in == 0) begin
					state<=5376;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=1487;
					out<=17;
				end
				if(in == 3) begin
					state<=7308;
					out<=18;
				end
				if(in == 4) begin
					state<=3419;
					out<=19;
				end
			end
			4356: begin
				if(in == 0) begin
					state<=5377;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=1488;
					out<=22;
				end
				if(in == 3) begin
					state<=7309;
					out<=23;
				end
				if(in == 4) begin
					state<=3420;
					out<=24;
				end
			end
			4357: begin
				if(in == 0) begin
					state<=5378;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=1489;
					out<=27;
				end
				if(in == 3) begin
					state<=7310;
					out<=28;
				end
				if(in == 4) begin
					state<=3421;
					out<=29;
				end
			end
			4358: begin
				if(in == 0) begin
					state<=5379;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=1490;
					out<=32;
				end
				if(in == 3) begin
					state<=7311;
					out<=33;
				end
				if(in == 4) begin
					state<=3422;
					out<=34;
				end
			end
			4359: begin
				if(in == 0) begin
					state<=5380;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=1491;
					out<=37;
				end
				if(in == 3) begin
					state<=7312;
					out<=38;
				end
				if(in == 4) begin
					state<=3423;
					out<=39;
				end
			end
			4360: begin
				if(in == 0) begin
					state<=5381;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=1492;
					out<=42;
				end
				if(in == 3) begin
					state<=7313;
					out<=43;
				end
				if(in == 4) begin
					state<=3424;
					out<=44;
				end
			end
			4361: begin
				if(in == 0) begin
					state<=5382;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=1493;
					out<=47;
				end
				if(in == 3) begin
					state<=7314;
					out<=48;
				end
				if(in == 4) begin
					state<=3425;
					out<=49;
				end
			end
			4362: begin
				if(in == 0) begin
					state<=5373;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=1484;
					out<=52;
				end
				if(in == 3) begin
					state<=7305;
					out<=53;
				end
				if(in == 4) begin
					state<=3416;
					out<=54;
				end
			end
			4363: begin
				if(in == 0) begin
					state<=4374;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=476;
					out<=57;
				end
				if(in == 3) begin
					state<=6363;
					out<=58;
				end
				if(in == 4) begin
					state<=2474;
					out<=59;
				end
			end
			4364: begin
				if(in == 0) begin
					state<=4375;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=477;
					out<=62;
				end
				if(in == 3) begin
					state<=6364;
					out<=63;
				end
				if(in == 4) begin
					state<=2475;
					out<=64;
				end
			end
			4365: begin
				if(in == 0) begin
					state<=4376;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=478;
					out<=67;
				end
				if(in == 3) begin
					state<=6365;
					out<=68;
				end
				if(in == 4) begin
					state<=2476;
					out<=69;
				end
			end
			4366: begin
				if(in == 0) begin
					state<=4377;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=479;
					out<=72;
				end
				if(in == 3) begin
					state<=6366;
					out<=73;
				end
				if(in == 4) begin
					state<=2477;
					out<=74;
				end
			end
			4367: begin
				if(in == 0) begin
					state<=4378;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=480;
					out<=77;
				end
				if(in == 3) begin
					state<=6367;
					out<=78;
				end
				if(in == 4) begin
					state<=2478;
					out<=79;
				end
			end
			4368: begin
				if(in == 0) begin
					state<=4379;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=481;
					out<=82;
				end
				if(in == 3) begin
					state<=6368;
					out<=83;
				end
				if(in == 4) begin
					state<=2479;
					out<=84;
				end
			end
			4369: begin
				if(in == 0) begin
					state<=4380;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=482;
					out<=87;
				end
				if(in == 3) begin
					state<=6369;
					out<=88;
				end
				if(in == 4) begin
					state<=2480;
					out<=89;
				end
			end
			4370: begin
				if(in == 0) begin
					state<=4381;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=483;
					out<=92;
				end
				if(in == 3) begin
					state<=6370;
					out<=93;
				end
				if(in == 4) begin
					state<=2481;
					out<=94;
				end
			end
			4371: begin
				if(in == 0) begin
					state<=4372;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=474;
					out<=97;
				end
				if(in == 3) begin
					state<=6361;
					out<=98;
				end
				if(in == 4) begin
					state<=2472;
					out<=99;
				end
			end
			4372: begin
				if(in == 0) begin
					state<=4383;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=485;
					out<=102;
				end
				if(in == 3) begin
					state<=6372;
					out<=103;
				end
				if(in == 4) begin
					state<=2483;
					out<=104;
				end
			end
			4373: begin
				if(in == 0) begin
					state<=4384;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=486;
					out<=107;
				end
				if(in == 3) begin
					state<=6373;
					out<=108;
				end
				if(in == 4) begin
					state<=2484;
					out<=109;
				end
			end
			4374: begin
				if(in == 0) begin
					state<=4385;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=487;
					out<=112;
				end
				if(in == 3) begin
					state<=6374;
					out<=113;
				end
				if(in == 4) begin
					state<=2485;
					out<=114;
				end
			end
			4375: begin
				if(in == 0) begin
					state<=4386;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=488;
					out<=117;
				end
				if(in == 3) begin
					state<=6375;
					out<=118;
				end
				if(in == 4) begin
					state<=2486;
					out<=119;
				end
			end
			4376: begin
				if(in == 0) begin
					state<=4387;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=489;
					out<=122;
				end
				if(in == 3) begin
					state<=6376;
					out<=123;
				end
				if(in == 4) begin
					state<=2487;
					out<=124;
				end
			end
			4377: begin
				if(in == 0) begin
					state<=4388;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=490;
					out<=127;
				end
				if(in == 3) begin
					state<=6377;
					out<=128;
				end
				if(in == 4) begin
					state<=2488;
					out<=129;
				end
			end
			4378: begin
				if(in == 0) begin
					state<=4389;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=491;
					out<=132;
				end
				if(in == 3) begin
					state<=6378;
					out<=133;
				end
				if(in == 4) begin
					state<=2489;
					out<=134;
				end
			end
			4379: begin
				if(in == 0) begin
					state<=4390;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=492;
					out<=137;
				end
				if(in == 3) begin
					state<=6379;
					out<=138;
				end
				if(in == 4) begin
					state<=2490;
					out<=139;
				end
			end
			4380: begin
				if(in == 0) begin
					state<=4391;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=493;
					out<=142;
				end
				if(in == 3) begin
					state<=6380;
					out<=143;
				end
				if(in == 4) begin
					state<=2491;
					out<=144;
				end
			end
			4381: begin
				if(in == 0) begin
					state<=4382;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=484;
					out<=147;
				end
				if(in == 3) begin
					state<=6371;
					out<=148;
				end
				if(in == 4) begin
					state<=2482;
					out<=149;
				end
			end
			4382: begin
				if(in == 0) begin
					state<=4393;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=495;
					out<=152;
				end
				if(in == 3) begin
					state<=6382;
					out<=153;
				end
				if(in == 4) begin
					state<=2493;
					out<=154;
				end
			end
			4383: begin
				if(in == 0) begin
					state<=4394;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=496;
					out<=157;
				end
				if(in == 3) begin
					state<=6383;
					out<=158;
				end
				if(in == 4) begin
					state<=2494;
					out<=159;
				end
			end
			4384: begin
				if(in == 0) begin
					state<=4395;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=497;
					out<=162;
				end
				if(in == 3) begin
					state<=6384;
					out<=163;
				end
				if(in == 4) begin
					state<=2495;
					out<=164;
				end
			end
			4385: begin
				if(in == 0) begin
					state<=4396;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=498;
					out<=167;
				end
				if(in == 3) begin
					state<=6385;
					out<=168;
				end
				if(in == 4) begin
					state<=2496;
					out<=169;
				end
			end
			4386: begin
				if(in == 0) begin
					state<=4397;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=499;
					out<=172;
				end
				if(in == 3) begin
					state<=6386;
					out<=173;
				end
				if(in == 4) begin
					state<=2497;
					out<=174;
				end
			end
			4387: begin
				if(in == 0) begin
					state<=4398;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=500;
					out<=177;
				end
				if(in == 3) begin
					state<=6387;
					out<=178;
				end
				if(in == 4) begin
					state<=2498;
					out<=179;
				end
			end
			4388: begin
				if(in == 0) begin
					state<=4399;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=501;
					out<=182;
				end
				if(in == 3) begin
					state<=6388;
					out<=183;
				end
				if(in == 4) begin
					state<=2499;
					out<=184;
				end
			end
			4389: begin
				if(in == 0) begin
					state<=4400;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=502;
					out<=187;
				end
				if(in == 3) begin
					state<=6389;
					out<=188;
				end
				if(in == 4) begin
					state<=2500;
					out<=189;
				end
			end
			4390: begin
				if(in == 0) begin
					state<=4401;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=503;
					out<=192;
				end
				if(in == 3) begin
					state<=6390;
					out<=193;
				end
				if(in == 4) begin
					state<=2501;
					out<=194;
				end
			end
			4391: begin
				if(in == 0) begin
					state<=4392;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=494;
					out<=197;
				end
				if(in == 3) begin
					state<=6381;
					out<=198;
				end
				if(in == 4) begin
					state<=2492;
					out<=199;
				end
			end
			4392: begin
				if(in == 0) begin
					state<=4403;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=505;
					out<=202;
				end
				if(in == 3) begin
					state<=6392;
					out<=203;
				end
				if(in == 4) begin
					state<=2503;
					out<=204;
				end
			end
			4393: begin
				if(in == 0) begin
					state<=4404;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=506;
					out<=207;
				end
				if(in == 3) begin
					state<=6393;
					out<=208;
				end
				if(in == 4) begin
					state<=2504;
					out<=209;
				end
			end
			4394: begin
				if(in == 0) begin
					state<=4405;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=507;
					out<=212;
				end
				if(in == 3) begin
					state<=6394;
					out<=213;
				end
				if(in == 4) begin
					state<=2505;
					out<=214;
				end
			end
			4395: begin
				if(in == 0) begin
					state<=4406;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=508;
					out<=217;
				end
				if(in == 3) begin
					state<=6395;
					out<=218;
				end
				if(in == 4) begin
					state<=2506;
					out<=219;
				end
			end
			4396: begin
				if(in == 0) begin
					state<=4407;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=509;
					out<=222;
				end
				if(in == 3) begin
					state<=6396;
					out<=223;
				end
				if(in == 4) begin
					state<=2507;
					out<=224;
				end
			end
			4397: begin
				if(in == 0) begin
					state<=4408;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=510;
					out<=227;
				end
				if(in == 3) begin
					state<=6397;
					out<=228;
				end
				if(in == 4) begin
					state<=2508;
					out<=229;
				end
			end
			4398: begin
				if(in == 0) begin
					state<=4409;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=511;
					out<=232;
				end
				if(in == 3) begin
					state<=6398;
					out<=233;
				end
				if(in == 4) begin
					state<=2509;
					out<=234;
				end
			end
			4399: begin
				if(in == 0) begin
					state<=4410;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=512;
					out<=237;
				end
				if(in == 3) begin
					state<=6399;
					out<=238;
				end
				if(in == 4) begin
					state<=2510;
					out<=239;
				end
			end
			4400: begin
				if(in == 0) begin
					state<=4411;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=513;
					out<=242;
				end
				if(in == 3) begin
					state<=6400;
					out<=243;
				end
				if(in == 4) begin
					state<=2511;
					out<=244;
				end
			end
			4401: begin
				if(in == 0) begin
					state<=4402;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=504;
					out<=247;
				end
				if(in == 3) begin
					state<=6391;
					out<=248;
				end
				if(in == 4) begin
					state<=2502;
					out<=249;
				end
			end
			4402: begin
				if(in == 0) begin
					state<=4413;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=515;
					out<=252;
				end
				if(in == 3) begin
					state<=6402;
					out<=253;
				end
				if(in == 4) begin
					state<=2513;
					out<=254;
				end
			end
			4403: begin
				if(in == 0) begin
					state<=4414;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=516;
					out<=1;
				end
				if(in == 3) begin
					state<=6403;
					out<=2;
				end
				if(in == 4) begin
					state<=2514;
					out<=3;
				end
			end
			4404: begin
				if(in == 0) begin
					state<=4415;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=517;
					out<=6;
				end
				if(in == 3) begin
					state<=6404;
					out<=7;
				end
				if(in == 4) begin
					state<=2515;
					out<=8;
				end
			end
			4405: begin
				if(in == 0) begin
					state<=4416;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=518;
					out<=11;
				end
				if(in == 3) begin
					state<=6405;
					out<=12;
				end
				if(in == 4) begin
					state<=2516;
					out<=13;
				end
			end
			4406: begin
				if(in == 0) begin
					state<=4417;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=519;
					out<=16;
				end
				if(in == 3) begin
					state<=6406;
					out<=17;
				end
				if(in == 4) begin
					state<=2517;
					out<=18;
				end
			end
			4407: begin
				if(in == 0) begin
					state<=4418;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=520;
					out<=21;
				end
				if(in == 3) begin
					state<=6407;
					out<=22;
				end
				if(in == 4) begin
					state<=2518;
					out<=23;
				end
			end
			4408: begin
				if(in == 0) begin
					state<=4419;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=521;
					out<=26;
				end
				if(in == 3) begin
					state<=6408;
					out<=27;
				end
				if(in == 4) begin
					state<=2519;
					out<=28;
				end
			end
			4409: begin
				if(in == 0) begin
					state<=4420;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=522;
					out<=31;
				end
				if(in == 3) begin
					state<=6409;
					out<=32;
				end
				if(in == 4) begin
					state<=2520;
					out<=33;
				end
			end
			4410: begin
				if(in == 0) begin
					state<=4421;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=523;
					out<=36;
				end
				if(in == 3) begin
					state<=6410;
					out<=37;
				end
				if(in == 4) begin
					state<=2521;
					out<=38;
				end
			end
			4411: begin
				if(in == 0) begin
					state<=4412;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=514;
					out<=41;
				end
				if(in == 3) begin
					state<=6401;
					out<=42;
				end
				if(in == 4) begin
					state<=2512;
					out<=43;
				end
			end
			4412: begin
				if(in == 0) begin
					state<=4423;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=525;
					out<=46;
				end
				if(in == 3) begin
					state<=6412;
					out<=47;
				end
				if(in == 4) begin
					state<=2523;
					out<=48;
				end
			end
			4413: begin
				if(in == 0) begin
					state<=4424;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=526;
					out<=51;
				end
				if(in == 3) begin
					state<=6413;
					out<=52;
				end
				if(in == 4) begin
					state<=2524;
					out<=53;
				end
			end
			4414: begin
				if(in == 0) begin
					state<=4425;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=527;
					out<=56;
				end
				if(in == 3) begin
					state<=6414;
					out<=57;
				end
				if(in == 4) begin
					state<=2525;
					out<=58;
				end
			end
			4415: begin
				if(in == 0) begin
					state<=4426;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=528;
					out<=61;
				end
				if(in == 3) begin
					state<=6415;
					out<=62;
				end
				if(in == 4) begin
					state<=2526;
					out<=63;
				end
			end
			4416: begin
				if(in == 0) begin
					state<=4427;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=529;
					out<=66;
				end
				if(in == 3) begin
					state<=6416;
					out<=67;
				end
				if(in == 4) begin
					state<=2527;
					out<=68;
				end
			end
			4417: begin
				if(in == 0) begin
					state<=4428;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=530;
					out<=71;
				end
				if(in == 3) begin
					state<=6417;
					out<=72;
				end
				if(in == 4) begin
					state<=2528;
					out<=73;
				end
			end
			4418: begin
				if(in == 0) begin
					state<=4429;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=531;
					out<=76;
				end
				if(in == 3) begin
					state<=6418;
					out<=77;
				end
				if(in == 4) begin
					state<=2529;
					out<=78;
				end
			end
			4419: begin
				if(in == 0) begin
					state<=4430;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=532;
					out<=81;
				end
				if(in == 3) begin
					state<=6419;
					out<=82;
				end
				if(in == 4) begin
					state<=2530;
					out<=83;
				end
			end
			4420: begin
				if(in == 0) begin
					state<=4431;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=533;
					out<=86;
				end
				if(in == 3) begin
					state<=6420;
					out<=87;
				end
				if(in == 4) begin
					state<=2531;
					out<=88;
				end
			end
			4421: begin
				if(in == 0) begin
					state<=4422;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=524;
					out<=91;
				end
				if(in == 3) begin
					state<=6411;
					out<=92;
				end
				if(in == 4) begin
					state<=2522;
					out<=93;
				end
			end
			4422: begin
				if(in == 0) begin
					state<=5405;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=1516;
					out<=96;
				end
				if(in == 3) begin
					state<=7337;
					out<=97;
				end
				if(in == 4) begin
					state<=3448;
					out<=98;
				end
			end
			4423: begin
				if(in == 0) begin
					state<=5406;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=1517;
					out<=101;
				end
				if(in == 3) begin
					state<=7338;
					out<=102;
				end
				if(in == 4) begin
					state<=3449;
					out<=103;
				end
			end
			4424: begin
				if(in == 0) begin
					state<=5407;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=1518;
					out<=106;
				end
				if(in == 3) begin
					state<=7339;
					out<=107;
				end
				if(in == 4) begin
					state<=3450;
					out<=108;
				end
			end
			4425: begin
				if(in == 0) begin
					state<=5408;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=1519;
					out<=111;
				end
				if(in == 3) begin
					state<=7340;
					out<=112;
				end
				if(in == 4) begin
					state<=3451;
					out<=113;
				end
			end
			4426: begin
				if(in == 0) begin
					state<=5409;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=1520;
					out<=116;
				end
				if(in == 3) begin
					state<=7341;
					out<=117;
				end
				if(in == 4) begin
					state<=3452;
					out<=118;
				end
			end
			4427: begin
				if(in == 0) begin
					state<=5410;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=1521;
					out<=121;
				end
				if(in == 3) begin
					state<=7342;
					out<=122;
				end
				if(in == 4) begin
					state<=3453;
					out<=123;
				end
			end
			4428: begin
				if(in == 0) begin
					state<=5411;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=1522;
					out<=126;
				end
				if(in == 3) begin
					state<=7343;
					out<=127;
				end
				if(in == 4) begin
					state<=3454;
					out<=128;
				end
			end
			4429: begin
				if(in == 0) begin
					state<=5412;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=1523;
					out<=131;
				end
				if(in == 3) begin
					state<=7344;
					out<=132;
				end
				if(in == 4) begin
					state<=3455;
					out<=133;
				end
			end
			4430: begin
				if(in == 0) begin
					state<=5413;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=1524;
					out<=136;
				end
				if(in == 3) begin
					state<=7345;
					out<=137;
				end
				if(in == 4) begin
					state<=3456;
					out<=138;
				end
			end
			4431: begin
				if(in == 0) begin
					state<=5404;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=1515;
					out<=141;
				end
				if(in == 3) begin
					state<=7336;
					out<=142;
				end
				if(in == 4) begin
					state<=3447;
					out<=143;
				end
			end
			4432: begin
				if(in == 0) begin
					state<=4443;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=545;
					out<=146;
				end
				if(in == 3) begin
					state<=6432;
					out<=147;
				end
				if(in == 4) begin
					state<=2543;
					out<=148;
				end
			end
			4433: begin
				if(in == 0) begin
					state<=4444;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=546;
					out<=151;
				end
				if(in == 3) begin
					state<=6433;
					out<=152;
				end
				if(in == 4) begin
					state<=2544;
					out<=153;
				end
			end
			4434: begin
				if(in == 0) begin
					state<=4445;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=547;
					out<=156;
				end
				if(in == 3) begin
					state<=6434;
					out<=157;
				end
				if(in == 4) begin
					state<=2545;
					out<=158;
				end
			end
			4435: begin
				if(in == 0) begin
					state<=4446;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=548;
					out<=161;
				end
				if(in == 3) begin
					state<=6435;
					out<=162;
				end
				if(in == 4) begin
					state<=2546;
					out<=163;
				end
			end
			4436: begin
				if(in == 0) begin
					state<=4447;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=549;
					out<=166;
				end
				if(in == 3) begin
					state<=6436;
					out<=167;
				end
				if(in == 4) begin
					state<=2547;
					out<=168;
				end
			end
			4437: begin
				if(in == 0) begin
					state<=4448;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=550;
					out<=171;
				end
				if(in == 3) begin
					state<=6437;
					out<=172;
				end
				if(in == 4) begin
					state<=2548;
					out<=173;
				end
			end
			4438: begin
				if(in == 0) begin
					state<=4449;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=551;
					out<=176;
				end
				if(in == 3) begin
					state<=6438;
					out<=177;
				end
				if(in == 4) begin
					state<=2549;
					out<=178;
				end
			end
			4439: begin
				if(in == 0) begin
					state<=4450;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=552;
					out<=181;
				end
				if(in == 3) begin
					state<=6439;
					out<=182;
				end
				if(in == 4) begin
					state<=2550;
					out<=183;
				end
			end
			4440: begin
				if(in == 0) begin
					state<=4441;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=543;
					out<=186;
				end
				if(in == 3) begin
					state<=6430;
					out<=187;
				end
				if(in == 4) begin
					state<=2541;
					out<=188;
				end
			end
			4441: begin
				if(in == 0) begin
					state<=4452;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=554;
					out<=191;
				end
				if(in == 3) begin
					state<=6441;
					out<=192;
				end
				if(in == 4) begin
					state<=2552;
					out<=193;
				end
			end
			4442: begin
				if(in == 0) begin
					state<=4453;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=555;
					out<=196;
				end
				if(in == 3) begin
					state<=6442;
					out<=197;
				end
				if(in == 4) begin
					state<=2553;
					out<=198;
				end
			end
			4443: begin
				if(in == 0) begin
					state<=4454;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=556;
					out<=201;
				end
				if(in == 3) begin
					state<=6443;
					out<=202;
				end
				if(in == 4) begin
					state<=2554;
					out<=203;
				end
			end
			4444: begin
				if(in == 0) begin
					state<=4455;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=557;
					out<=206;
				end
				if(in == 3) begin
					state<=6444;
					out<=207;
				end
				if(in == 4) begin
					state<=2555;
					out<=208;
				end
			end
			4445: begin
				if(in == 0) begin
					state<=4456;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=558;
					out<=211;
				end
				if(in == 3) begin
					state<=6445;
					out<=212;
				end
				if(in == 4) begin
					state<=2556;
					out<=213;
				end
			end
			4446: begin
				if(in == 0) begin
					state<=4457;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=559;
					out<=216;
				end
				if(in == 3) begin
					state<=6446;
					out<=217;
				end
				if(in == 4) begin
					state<=2557;
					out<=218;
				end
			end
			4447: begin
				if(in == 0) begin
					state<=4458;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=560;
					out<=221;
				end
				if(in == 3) begin
					state<=6447;
					out<=222;
				end
				if(in == 4) begin
					state<=2558;
					out<=223;
				end
			end
			4448: begin
				if(in == 0) begin
					state<=4459;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=561;
					out<=226;
				end
				if(in == 3) begin
					state<=6448;
					out<=227;
				end
				if(in == 4) begin
					state<=2559;
					out<=228;
				end
			end
			4449: begin
				if(in == 0) begin
					state<=4460;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=562;
					out<=231;
				end
				if(in == 3) begin
					state<=6449;
					out<=232;
				end
				if(in == 4) begin
					state<=2560;
					out<=233;
				end
			end
			4450: begin
				if(in == 0) begin
					state<=4451;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=553;
					out<=236;
				end
				if(in == 3) begin
					state<=6440;
					out<=237;
				end
				if(in == 4) begin
					state<=2551;
					out<=238;
				end
			end
			4451: begin
				if(in == 0) begin
					state<=4462;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=564;
					out<=241;
				end
				if(in == 3) begin
					state<=6451;
					out<=242;
				end
				if(in == 4) begin
					state<=2562;
					out<=243;
				end
			end
			4452: begin
				if(in == 0) begin
					state<=4463;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=565;
					out<=246;
				end
				if(in == 3) begin
					state<=6452;
					out<=247;
				end
				if(in == 4) begin
					state<=2563;
					out<=248;
				end
			end
			4453: begin
				if(in == 0) begin
					state<=4464;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=566;
					out<=251;
				end
				if(in == 3) begin
					state<=6453;
					out<=252;
				end
				if(in == 4) begin
					state<=2564;
					out<=253;
				end
			end
			4454: begin
				if(in == 0) begin
					state<=4465;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=567;
					out<=0;
				end
				if(in == 3) begin
					state<=6454;
					out<=1;
				end
				if(in == 4) begin
					state<=2565;
					out<=2;
				end
			end
			4455: begin
				if(in == 0) begin
					state<=4466;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=568;
					out<=5;
				end
				if(in == 3) begin
					state<=6455;
					out<=6;
				end
				if(in == 4) begin
					state<=2566;
					out<=7;
				end
			end
			4456: begin
				if(in == 0) begin
					state<=4467;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=569;
					out<=10;
				end
				if(in == 3) begin
					state<=6456;
					out<=11;
				end
				if(in == 4) begin
					state<=2567;
					out<=12;
				end
			end
			4457: begin
				if(in == 0) begin
					state<=4468;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=570;
					out<=15;
				end
				if(in == 3) begin
					state<=6457;
					out<=16;
				end
				if(in == 4) begin
					state<=2568;
					out<=17;
				end
			end
			4458: begin
				if(in == 0) begin
					state<=4469;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=571;
					out<=20;
				end
				if(in == 3) begin
					state<=6458;
					out<=21;
				end
				if(in == 4) begin
					state<=2569;
					out<=22;
				end
			end
			4459: begin
				if(in == 0) begin
					state<=4470;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=572;
					out<=25;
				end
				if(in == 3) begin
					state<=6459;
					out<=26;
				end
				if(in == 4) begin
					state<=2570;
					out<=27;
				end
			end
			4460: begin
				if(in == 0) begin
					state<=4461;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=563;
					out<=30;
				end
				if(in == 3) begin
					state<=6450;
					out<=31;
				end
				if(in == 4) begin
					state<=2561;
					out<=32;
				end
			end
			4461: begin
				if(in == 0) begin
					state<=4472;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=574;
					out<=35;
				end
				if(in == 3) begin
					state<=6461;
					out<=36;
				end
				if(in == 4) begin
					state<=2572;
					out<=37;
				end
			end
			4462: begin
				if(in == 0) begin
					state<=4473;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=575;
					out<=40;
				end
				if(in == 3) begin
					state<=6462;
					out<=41;
				end
				if(in == 4) begin
					state<=2573;
					out<=42;
				end
			end
			4463: begin
				if(in == 0) begin
					state<=4474;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=576;
					out<=45;
				end
				if(in == 3) begin
					state<=6463;
					out<=46;
				end
				if(in == 4) begin
					state<=2574;
					out<=47;
				end
			end
			4464: begin
				if(in == 0) begin
					state<=4475;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=577;
					out<=50;
				end
				if(in == 3) begin
					state<=6464;
					out<=51;
				end
				if(in == 4) begin
					state<=2575;
					out<=52;
				end
			end
			4465: begin
				if(in == 0) begin
					state<=4476;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=578;
					out<=55;
				end
				if(in == 3) begin
					state<=6465;
					out<=56;
				end
				if(in == 4) begin
					state<=2576;
					out<=57;
				end
			end
			4466: begin
				if(in == 0) begin
					state<=4477;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=579;
					out<=60;
				end
				if(in == 3) begin
					state<=6466;
					out<=61;
				end
				if(in == 4) begin
					state<=2577;
					out<=62;
				end
			end
			4467: begin
				if(in == 0) begin
					state<=4478;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=580;
					out<=65;
				end
				if(in == 3) begin
					state<=6467;
					out<=66;
				end
				if(in == 4) begin
					state<=2578;
					out<=67;
				end
			end
			4468: begin
				if(in == 0) begin
					state<=4479;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=581;
					out<=70;
				end
				if(in == 3) begin
					state<=6468;
					out<=71;
				end
				if(in == 4) begin
					state<=2579;
					out<=72;
				end
			end
			4469: begin
				if(in == 0) begin
					state<=4480;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=582;
					out<=75;
				end
				if(in == 3) begin
					state<=6469;
					out<=76;
				end
				if(in == 4) begin
					state<=2580;
					out<=77;
				end
			end
			4470: begin
				if(in == 0) begin
					state<=4471;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=573;
					out<=80;
				end
				if(in == 3) begin
					state<=6460;
					out<=81;
				end
				if(in == 4) begin
					state<=2571;
					out<=82;
				end
			end
			4471: begin
				if(in == 0) begin
					state<=4482;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=584;
					out<=85;
				end
				if(in == 3) begin
					state<=6471;
					out<=86;
				end
				if(in == 4) begin
					state<=2582;
					out<=87;
				end
			end
			4472: begin
				if(in == 0) begin
					state<=4483;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=585;
					out<=90;
				end
				if(in == 3) begin
					state<=6472;
					out<=91;
				end
				if(in == 4) begin
					state<=2583;
					out<=92;
				end
			end
			4473: begin
				if(in == 0) begin
					state<=4484;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=586;
					out<=95;
				end
				if(in == 3) begin
					state<=6473;
					out<=96;
				end
				if(in == 4) begin
					state<=2584;
					out<=97;
				end
			end
			4474: begin
				if(in == 0) begin
					state<=4485;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=587;
					out<=100;
				end
				if(in == 3) begin
					state<=6474;
					out<=101;
				end
				if(in == 4) begin
					state<=2585;
					out<=102;
				end
			end
			4475: begin
				if(in == 0) begin
					state<=4486;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=588;
					out<=105;
				end
				if(in == 3) begin
					state<=6475;
					out<=106;
				end
				if(in == 4) begin
					state<=2586;
					out<=107;
				end
			end
			4476: begin
				if(in == 0) begin
					state<=4487;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=589;
					out<=110;
				end
				if(in == 3) begin
					state<=6476;
					out<=111;
				end
				if(in == 4) begin
					state<=2587;
					out<=112;
				end
			end
			4477: begin
				if(in == 0) begin
					state<=4488;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=590;
					out<=115;
				end
				if(in == 3) begin
					state<=6477;
					out<=116;
				end
				if(in == 4) begin
					state<=2588;
					out<=117;
				end
			end
			4478: begin
				if(in == 0) begin
					state<=4489;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=591;
					out<=120;
				end
				if(in == 3) begin
					state<=6478;
					out<=121;
				end
				if(in == 4) begin
					state<=2589;
					out<=122;
				end
			end
			4479: begin
				if(in == 0) begin
					state<=4490;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=592;
					out<=125;
				end
				if(in == 3) begin
					state<=6479;
					out<=126;
				end
				if(in == 4) begin
					state<=2590;
					out<=127;
				end
			end
			4480: begin
				if(in == 0) begin
					state<=4481;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=583;
					out<=130;
				end
				if(in == 3) begin
					state<=6470;
					out<=131;
				end
				if(in == 4) begin
					state<=2581;
					out<=132;
				end
			end
			4481: begin
				if(in == 0) begin
					state<=4492;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=594;
					out<=135;
				end
				if(in == 3) begin
					state<=6481;
					out<=136;
				end
				if(in == 4) begin
					state<=2592;
					out<=137;
				end
			end
			4482: begin
				if(in == 0) begin
					state<=4493;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=595;
					out<=140;
				end
				if(in == 3) begin
					state<=6482;
					out<=141;
				end
				if(in == 4) begin
					state<=2593;
					out<=142;
				end
			end
			4483: begin
				if(in == 0) begin
					state<=4494;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=596;
					out<=145;
				end
				if(in == 3) begin
					state<=6483;
					out<=146;
				end
				if(in == 4) begin
					state<=2594;
					out<=147;
				end
			end
			4484: begin
				if(in == 0) begin
					state<=4495;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=597;
					out<=150;
				end
				if(in == 3) begin
					state<=6484;
					out<=151;
				end
				if(in == 4) begin
					state<=2595;
					out<=152;
				end
			end
			4485: begin
				if(in == 0) begin
					state<=4496;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=598;
					out<=155;
				end
				if(in == 3) begin
					state<=6485;
					out<=156;
				end
				if(in == 4) begin
					state<=2596;
					out<=157;
				end
			end
			4486: begin
				if(in == 0) begin
					state<=4497;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=599;
					out<=160;
				end
				if(in == 3) begin
					state<=6486;
					out<=161;
				end
				if(in == 4) begin
					state<=2597;
					out<=162;
				end
			end
			4487: begin
				if(in == 0) begin
					state<=4498;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=600;
					out<=165;
				end
				if(in == 3) begin
					state<=6487;
					out<=166;
				end
				if(in == 4) begin
					state<=2598;
					out<=167;
				end
			end
			4488: begin
				if(in == 0) begin
					state<=4499;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=601;
					out<=170;
				end
				if(in == 3) begin
					state<=6488;
					out<=171;
				end
				if(in == 4) begin
					state<=2599;
					out<=172;
				end
			end
			4489: begin
				if(in == 0) begin
					state<=4500;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=602;
					out<=175;
				end
				if(in == 3) begin
					state<=6489;
					out<=176;
				end
				if(in == 4) begin
					state<=2600;
					out<=177;
				end
			end
			4490: begin
				if(in == 0) begin
					state<=4491;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=593;
					out<=180;
				end
				if(in == 3) begin
					state<=6480;
					out<=181;
				end
				if(in == 4) begin
					state<=2591;
					out<=182;
				end
			end
			4491: begin
				if(in == 0) begin
					state<=5436;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=1547;
					out<=185;
				end
				if(in == 3) begin
					state<=7368;
					out<=186;
				end
				if(in == 4) begin
					state<=3479;
					out<=187;
				end
			end
			4492: begin
				if(in == 0) begin
					state<=5437;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=1548;
					out<=190;
				end
				if(in == 3) begin
					state<=7369;
					out<=191;
				end
				if(in == 4) begin
					state<=3480;
					out<=192;
				end
			end
			4493: begin
				if(in == 0) begin
					state<=5438;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=1549;
					out<=195;
				end
				if(in == 3) begin
					state<=7370;
					out<=196;
				end
				if(in == 4) begin
					state<=3481;
					out<=197;
				end
			end
			4494: begin
				if(in == 0) begin
					state<=5439;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=1550;
					out<=200;
				end
				if(in == 3) begin
					state<=7371;
					out<=201;
				end
				if(in == 4) begin
					state<=3482;
					out<=202;
				end
			end
			4495: begin
				if(in == 0) begin
					state<=5440;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=1551;
					out<=205;
				end
				if(in == 3) begin
					state<=7372;
					out<=206;
				end
				if(in == 4) begin
					state<=3483;
					out<=207;
				end
			end
			4496: begin
				if(in == 0) begin
					state<=5441;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=1552;
					out<=210;
				end
				if(in == 3) begin
					state<=7373;
					out<=211;
				end
				if(in == 4) begin
					state<=3484;
					out<=212;
				end
			end
			4497: begin
				if(in == 0) begin
					state<=5442;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=1553;
					out<=215;
				end
				if(in == 3) begin
					state<=7374;
					out<=216;
				end
				if(in == 4) begin
					state<=3485;
					out<=217;
				end
			end
			4498: begin
				if(in == 0) begin
					state<=5443;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=1554;
					out<=220;
				end
				if(in == 3) begin
					state<=7375;
					out<=221;
				end
				if(in == 4) begin
					state<=3486;
					out<=222;
				end
			end
			4499: begin
				if(in == 0) begin
					state<=5444;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=1555;
					out<=225;
				end
				if(in == 3) begin
					state<=7376;
					out<=226;
				end
				if(in == 4) begin
					state<=3487;
					out<=227;
				end
			end
			4500: begin
				if(in == 0) begin
					state<=5435;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=1546;
					out<=230;
				end
				if(in == 3) begin
					state<=7367;
					out<=231;
				end
				if(in == 4) begin
					state<=3478;
					out<=232;
				end
			end
			4501: begin
				if(in == 0) begin
					state<=4512;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=614;
					out<=235;
				end
				if(in == 3) begin
					state<=6501;
					out<=236;
				end
				if(in == 4) begin
					state<=2612;
					out<=237;
				end
			end
			4502: begin
				if(in == 0) begin
					state<=4513;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=615;
					out<=240;
				end
				if(in == 3) begin
					state<=6502;
					out<=241;
				end
				if(in == 4) begin
					state<=2613;
					out<=242;
				end
			end
			4503: begin
				if(in == 0) begin
					state<=4514;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=616;
					out<=245;
				end
				if(in == 3) begin
					state<=6503;
					out<=246;
				end
				if(in == 4) begin
					state<=2614;
					out<=247;
				end
			end
			4504: begin
				if(in == 0) begin
					state<=4515;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=617;
					out<=250;
				end
				if(in == 3) begin
					state<=6504;
					out<=251;
				end
				if(in == 4) begin
					state<=2615;
					out<=252;
				end
			end
			4505: begin
				if(in == 0) begin
					state<=4516;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=618;
					out<=255;
				end
				if(in == 3) begin
					state<=6505;
					out<=0;
				end
				if(in == 4) begin
					state<=2616;
					out<=1;
				end
			end
			4506: begin
				if(in == 0) begin
					state<=4517;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=619;
					out<=4;
				end
				if(in == 3) begin
					state<=6506;
					out<=5;
				end
				if(in == 4) begin
					state<=2617;
					out<=6;
				end
			end
			4507: begin
				if(in == 0) begin
					state<=4518;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=620;
					out<=9;
				end
				if(in == 3) begin
					state<=6507;
					out<=10;
				end
				if(in == 4) begin
					state<=2618;
					out<=11;
				end
			end
			4508: begin
				if(in == 0) begin
					state<=4519;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=621;
					out<=14;
				end
				if(in == 3) begin
					state<=6508;
					out<=15;
				end
				if(in == 4) begin
					state<=2619;
					out<=16;
				end
			end
			4509: begin
				if(in == 0) begin
					state<=4510;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=612;
					out<=19;
				end
				if(in == 3) begin
					state<=6499;
					out<=20;
				end
				if(in == 4) begin
					state<=2610;
					out<=21;
				end
			end
			4510: begin
				if(in == 0) begin
					state<=4521;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=623;
					out<=24;
				end
				if(in == 3) begin
					state<=6510;
					out<=25;
				end
				if(in == 4) begin
					state<=2621;
					out<=26;
				end
			end
			4511: begin
				if(in == 0) begin
					state<=4522;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=624;
					out<=29;
				end
				if(in == 3) begin
					state<=6511;
					out<=30;
				end
				if(in == 4) begin
					state<=2622;
					out<=31;
				end
			end
			4512: begin
				if(in == 0) begin
					state<=4523;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=625;
					out<=34;
				end
				if(in == 3) begin
					state<=6512;
					out<=35;
				end
				if(in == 4) begin
					state<=2623;
					out<=36;
				end
			end
			4513: begin
				if(in == 0) begin
					state<=4524;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=626;
					out<=39;
				end
				if(in == 3) begin
					state<=6513;
					out<=40;
				end
				if(in == 4) begin
					state<=2624;
					out<=41;
				end
			end
			4514: begin
				if(in == 0) begin
					state<=4525;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=627;
					out<=44;
				end
				if(in == 3) begin
					state<=6514;
					out<=45;
				end
				if(in == 4) begin
					state<=2625;
					out<=46;
				end
			end
			4515: begin
				if(in == 0) begin
					state<=4526;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=628;
					out<=49;
				end
				if(in == 3) begin
					state<=6515;
					out<=50;
				end
				if(in == 4) begin
					state<=2626;
					out<=51;
				end
			end
			4516: begin
				if(in == 0) begin
					state<=4527;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=629;
					out<=54;
				end
				if(in == 3) begin
					state<=6516;
					out<=55;
				end
				if(in == 4) begin
					state<=2627;
					out<=56;
				end
			end
			4517: begin
				if(in == 0) begin
					state<=4528;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=630;
					out<=59;
				end
				if(in == 3) begin
					state<=6517;
					out<=60;
				end
				if(in == 4) begin
					state<=2628;
					out<=61;
				end
			end
			4518: begin
				if(in == 0) begin
					state<=4529;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=631;
					out<=64;
				end
				if(in == 3) begin
					state<=6518;
					out<=65;
				end
				if(in == 4) begin
					state<=2629;
					out<=66;
				end
			end
			4519: begin
				if(in == 0) begin
					state<=4520;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=622;
					out<=69;
				end
				if(in == 3) begin
					state<=6509;
					out<=70;
				end
				if(in == 4) begin
					state<=2620;
					out<=71;
				end
			end
			4520: begin
				if(in == 0) begin
					state<=4531;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=633;
					out<=74;
				end
				if(in == 3) begin
					state<=6520;
					out<=75;
				end
				if(in == 4) begin
					state<=2631;
					out<=76;
				end
			end
			4521: begin
				if(in == 0) begin
					state<=4532;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=634;
					out<=79;
				end
				if(in == 3) begin
					state<=6521;
					out<=80;
				end
				if(in == 4) begin
					state<=2632;
					out<=81;
				end
			end
			4522: begin
				if(in == 0) begin
					state<=4533;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=635;
					out<=84;
				end
				if(in == 3) begin
					state<=6522;
					out<=85;
				end
				if(in == 4) begin
					state<=2633;
					out<=86;
				end
			end
			4523: begin
				if(in == 0) begin
					state<=4534;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=636;
					out<=89;
				end
				if(in == 3) begin
					state<=6523;
					out<=90;
				end
				if(in == 4) begin
					state<=2634;
					out<=91;
				end
			end
			4524: begin
				if(in == 0) begin
					state<=4535;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=637;
					out<=94;
				end
				if(in == 3) begin
					state<=6524;
					out<=95;
				end
				if(in == 4) begin
					state<=2635;
					out<=96;
				end
			end
			4525: begin
				if(in == 0) begin
					state<=4536;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=638;
					out<=99;
				end
				if(in == 3) begin
					state<=6525;
					out<=100;
				end
				if(in == 4) begin
					state<=2636;
					out<=101;
				end
			end
			4526: begin
				if(in == 0) begin
					state<=4537;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=639;
					out<=104;
				end
				if(in == 3) begin
					state<=6526;
					out<=105;
				end
				if(in == 4) begin
					state<=2637;
					out<=106;
				end
			end
			4527: begin
				if(in == 0) begin
					state<=4538;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=640;
					out<=109;
				end
				if(in == 3) begin
					state<=6527;
					out<=110;
				end
				if(in == 4) begin
					state<=2638;
					out<=111;
				end
			end
			4528: begin
				if(in == 0) begin
					state<=4539;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=641;
					out<=114;
				end
				if(in == 3) begin
					state<=6528;
					out<=115;
				end
				if(in == 4) begin
					state<=2639;
					out<=116;
				end
			end
			4529: begin
				if(in == 0) begin
					state<=4530;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=632;
					out<=119;
				end
				if(in == 3) begin
					state<=6519;
					out<=120;
				end
				if(in == 4) begin
					state<=2630;
					out<=121;
				end
			end
			4530: begin
				if(in == 0) begin
					state<=4541;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=643;
					out<=124;
				end
				if(in == 3) begin
					state<=6530;
					out<=125;
				end
				if(in == 4) begin
					state<=2641;
					out<=126;
				end
			end
			4531: begin
				if(in == 0) begin
					state<=4542;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=644;
					out<=129;
				end
				if(in == 3) begin
					state<=6531;
					out<=130;
				end
				if(in == 4) begin
					state<=2642;
					out<=131;
				end
			end
			4532: begin
				if(in == 0) begin
					state<=4543;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=645;
					out<=134;
				end
				if(in == 3) begin
					state<=6532;
					out<=135;
				end
				if(in == 4) begin
					state<=2643;
					out<=136;
				end
			end
			4533: begin
				if(in == 0) begin
					state<=4544;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=646;
					out<=139;
				end
				if(in == 3) begin
					state<=6533;
					out<=140;
				end
				if(in == 4) begin
					state<=2644;
					out<=141;
				end
			end
			4534: begin
				if(in == 0) begin
					state<=4545;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=647;
					out<=144;
				end
				if(in == 3) begin
					state<=6534;
					out<=145;
				end
				if(in == 4) begin
					state<=2645;
					out<=146;
				end
			end
			4535: begin
				if(in == 0) begin
					state<=4546;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=648;
					out<=149;
				end
				if(in == 3) begin
					state<=6535;
					out<=150;
				end
				if(in == 4) begin
					state<=2646;
					out<=151;
				end
			end
			4536: begin
				if(in == 0) begin
					state<=4547;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=649;
					out<=154;
				end
				if(in == 3) begin
					state<=6536;
					out<=155;
				end
				if(in == 4) begin
					state<=2647;
					out<=156;
				end
			end
			4537: begin
				if(in == 0) begin
					state<=4548;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=650;
					out<=159;
				end
				if(in == 3) begin
					state<=6537;
					out<=160;
				end
				if(in == 4) begin
					state<=2648;
					out<=161;
				end
			end
			4538: begin
				if(in == 0) begin
					state<=4549;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=651;
					out<=164;
				end
				if(in == 3) begin
					state<=6538;
					out<=165;
				end
				if(in == 4) begin
					state<=2649;
					out<=166;
				end
			end
			4539: begin
				if(in == 0) begin
					state<=4540;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=642;
					out<=169;
				end
				if(in == 3) begin
					state<=6529;
					out<=170;
				end
				if(in == 4) begin
					state<=2640;
					out<=171;
				end
			end
			4540: begin
				if(in == 0) begin
					state<=4551;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=653;
					out<=174;
				end
				if(in == 3) begin
					state<=6540;
					out<=175;
				end
				if(in == 4) begin
					state<=2651;
					out<=176;
				end
			end
			4541: begin
				if(in == 0) begin
					state<=4552;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=654;
					out<=179;
				end
				if(in == 3) begin
					state<=6541;
					out<=180;
				end
				if(in == 4) begin
					state<=2652;
					out<=181;
				end
			end
			4542: begin
				if(in == 0) begin
					state<=4553;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=655;
					out<=184;
				end
				if(in == 3) begin
					state<=6542;
					out<=185;
				end
				if(in == 4) begin
					state<=2653;
					out<=186;
				end
			end
			4543: begin
				if(in == 0) begin
					state<=4554;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=656;
					out<=189;
				end
				if(in == 3) begin
					state<=6543;
					out<=190;
				end
				if(in == 4) begin
					state<=2654;
					out<=191;
				end
			end
			4544: begin
				if(in == 0) begin
					state<=4555;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=657;
					out<=194;
				end
				if(in == 3) begin
					state<=6544;
					out<=195;
				end
				if(in == 4) begin
					state<=2655;
					out<=196;
				end
			end
			4545: begin
				if(in == 0) begin
					state<=4556;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=658;
					out<=199;
				end
				if(in == 3) begin
					state<=6545;
					out<=200;
				end
				if(in == 4) begin
					state<=2656;
					out<=201;
				end
			end
			4546: begin
				if(in == 0) begin
					state<=4557;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=659;
					out<=204;
				end
				if(in == 3) begin
					state<=6546;
					out<=205;
				end
				if(in == 4) begin
					state<=2657;
					out<=206;
				end
			end
			4547: begin
				if(in == 0) begin
					state<=4558;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=660;
					out<=209;
				end
				if(in == 3) begin
					state<=6547;
					out<=210;
				end
				if(in == 4) begin
					state<=2658;
					out<=211;
				end
			end
			4548: begin
				if(in == 0) begin
					state<=4559;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=661;
					out<=214;
				end
				if(in == 3) begin
					state<=6548;
					out<=215;
				end
				if(in == 4) begin
					state<=2659;
					out<=216;
				end
			end
			4549: begin
				if(in == 0) begin
					state<=4550;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=652;
					out<=219;
				end
				if(in == 3) begin
					state<=6539;
					out<=220;
				end
				if(in == 4) begin
					state<=2650;
					out<=221;
				end
			end
			4550: begin
				if(in == 0) begin
					state<=4561;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=663;
					out<=224;
				end
				if(in == 3) begin
					state<=6550;
					out<=225;
				end
				if(in == 4) begin
					state<=2661;
					out<=226;
				end
			end
			4551: begin
				if(in == 0) begin
					state<=4562;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=664;
					out<=229;
				end
				if(in == 3) begin
					state<=6551;
					out<=230;
				end
				if(in == 4) begin
					state<=2662;
					out<=231;
				end
			end
			4552: begin
				if(in == 0) begin
					state<=4563;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=665;
					out<=234;
				end
				if(in == 3) begin
					state<=6552;
					out<=235;
				end
				if(in == 4) begin
					state<=2663;
					out<=236;
				end
			end
			4553: begin
				if(in == 0) begin
					state<=4564;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=666;
					out<=239;
				end
				if(in == 3) begin
					state<=6553;
					out<=240;
				end
				if(in == 4) begin
					state<=2664;
					out<=241;
				end
			end
			4554: begin
				if(in == 0) begin
					state<=4565;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=667;
					out<=244;
				end
				if(in == 3) begin
					state<=6554;
					out<=245;
				end
				if(in == 4) begin
					state<=2665;
					out<=246;
				end
			end
			4555: begin
				if(in == 0) begin
					state<=4566;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=668;
					out<=249;
				end
				if(in == 3) begin
					state<=6555;
					out<=250;
				end
				if(in == 4) begin
					state<=2666;
					out<=251;
				end
			end
			4556: begin
				if(in == 0) begin
					state<=4567;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=669;
					out<=254;
				end
				if(in == 3) begin
					state<=6556;
					out<=255;
				end
				if(in == 4) begin
					state<=2667;
					out<=0;
				end
			end
			4557: begin
				if(in == 0) begin
					state<=4568;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=670;
					out<=3;
				end
				if(in == 3) begin
					state<=6557;
					out<=4;
				end
				if(in == 4) begin
					state<=2668;
					out<=5;
				end
			end
			4558: begin
				if(in == 0) begin
					state<=4569;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=671;
					out<=8;
				end
				if(in == 3) begin
					state<=6558;
					out<=9;
				end
				if(in == 4) begin
					state<=2669;
					out<=10;
				end
			end
			4559: begin
				if(in == 0) begin
					state<=4560;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=662;
					out<=13;
				end
				if(in == 3) begin
					state<=6549;
					out<=14;
				end
				if(in == 4) begin
					state<=2660;
					out<=15;
				end
			end
			4560: begin
				if(in == 0) begin
					state<=5467;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=1578;
					out<=18;
				end
				if(in == 3) begin
					state<=7120;
					out<=19;
				end
				if(in == 4) begin
					state<=3231;
					out<=20;
				end
			end
			4561: begin
				if(in == 0) begin
					state<=5468;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=1579;
					out<=23;
				end
				if(in == 3) begin
					state<=7121;
					out<=24;
				end
				if(in == 4) begin
					state<=3232;
					out<=25;
				end
			end
			4562: begin
				if(in == 0) begin
					state<=5469;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=1580;
					out<=28;
				end
				if(in == 3) begin
					state<=7122;
					out<=29;
				end
				if(in == 4) begin
					state<=3233;
					out<=30;
				end
			end
			4563: begin
				if(in == 0) begin
					state<=5470;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=1581;
					out<=33;
				end
				if(in == 3) begin
					state<=7123;
					out<=34;
				end
				if(in == 4) begin
					state<=3234;
					out<=35;
				end
			end
			4564: begin
				if(in == 0) begin
					state<=5471;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=1582;
					out<=38;
				end
				if(in == 3) begin
					state<=7124;
					out<=39;
				end
				if(in == 4) begin
					state<=3235;
					out<=40;
				end
			end
			4565: begin
				if(in == 0) begin
					state<=5472;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=1583;
					out<=43;
				end
				if(in == 3) begin
					state<=7125;
					out<=44;
				end
				if(in == 4) begin
					state<=3236;
					out<=45;
				end
			end
			4566: begin
				if(in == 0) begin
					state<=5473;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=1584;
					out<=48;
				end
				if(in == 3) begin
					state<=7126;
					out<=49;
				end
				if(in == 4) begin
					state<=3237;
					out<=50;
				end
			end
			4567: begin
				if(in == 0) begin
					state<=5474;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=1585;
					out<=53;
				end
				if(in == 3) begin
					state<=7127;
					out<=54;
				end
				if(in == 4) begin
					state<=3238;
					out<=55;
				end
			end
			4568: begin
				if(in == 0) begin
					state<=5475;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=1586;
					out<=58;
				end
				if(in == 3) begin
					state<=7128;
					out<=59;
				end
				if(in == 4) begin
					state<=3239;
					out<=60;
				end
			end
			4569: begin
				if(in == 0) begin
					state<=5466;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=1577;
					out<=63;
				end
				if(in == 3) begin
					state<=7119;
					out<=64;
				end
				if(in == 4) begin
					state<=3230;
					out<=65;
				end
			end
			4570: begin
				if(in == 0) begin
					state<=4581;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=683;
					out<=68;
				end
				if(in == 3) begin
					state<=6570;
					out<=69;
				end
				if(in == 4) begin
					state<=2681;
					out<=70;
				end
			end
			4571: begin
				if(in == 0) begin
					state<=4582;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=684;
					out<=73;
				end
				if(in == 3) begin
					state<=6571;
					out<=74;
				end
				if(in == 4) begin
					state<=2682;
					out<=75;
				end
			end
			4572: begin
				if(in == 0) begin
					state<=4583;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=685;
					out<=78;
				end
				if(in == 3) begin
					state<=6572;
					out<=79;
				end
				if(in == 4) begin
					state<=2683;
					out<=80;
				end
			end
			4573: begin
				if(in == 0) begin
					state<=4584;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=686;
					out<=83;
				end
				if(in == 3) begin
					state<=6573;
					out<=84;
				end
				if(in == 4) begin
					state<=2684;
					out<=85;
				end
			end
			4574: begin
				if(in == 0) begin
					state<=4585;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=687;
					out<=88;
				end
				if(in == 3) begin
					state<=6574;
					out<=89;
				end
				if(in == 4) begin
					state<=2685;
					out<=90;
				end
			end
			4575: begin
				if(in == 0) begin
					state<=4586;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=688;
					out<=93;
				end
				if(in == 3) begin
					state<=6575;
					out<=94;
				end
				if(in == 4) begin
					state<=2686;
					out<=95;
				end
			end
			4576: begin
				if(in == 0) begin
					state<=4587;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=689;
					out<=98;
				end
				if(in == 3) begin
					state<=6576;
					out<=99;
				end
				if(in == 4) begin
					state<=2687;
					out<=100;
				end
			end
			4577: begin
				if(in == 0) begin
					state<=4588;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=690;
					out<=103;
				end
				if(in == 3) begin
					state<=6577;
					out<=104;
				end
				if(in == 4) begin
					state<=2688;
					out<=105;
				end
			end
			4578: begin
				if(in == 0) begin
					state<=4579;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=681;
					out<=108;
				end
				if(in == 3) begin
					state<=6568;
					out<=109;
				end
				if(in == 4) begin
					state<=2679;
					out<=110;
				end
			end
			4579: begin
				if(in == 0) begin
					state<=3900;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=2;
					out<=113;
				end
				if(in == 3) begin
					state<=5889;
					out<=114;
				end
				if(in == 4) begin
					state<=2000;
					out<=115;
				end
			end
			4580: begin
				if(in == 0) begin
					state<=3901;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=3;
					out<=118;
				end
				if(in == 3) begin
					state<=5890;
					out<=119;
				end
				if(in == 4) begin
					state<=2001;
					out<=120;
				end
			end
			4581: begin
				if(in == 0) begin
					state<=3902;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=4;
					out<=123;
				end
				if(in == 3) begin
					state<=5891;
					out<=124;
				end
				if(in == 4) begin
					state<=2002;
					out<=125;
				end
			end
			4582: begin
				if(in == 0) begin
					state<=3903;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=5;
					out<=128;
				end
				if(in == 3) begin
					state<=5892;
					out<=129;
				end
				if(in == 4) begin
					state<=2003;
					out<=130;
				end
			end
			4583: begin
				if(in == 0) begin
					state<=3904;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=6;
					out<=133;
				end
				if(in == 3) begin
					state<=5893;
					out<=134;
				end
				if(in == 4) begin
					state<=2004;
					out<=135;
				end
			end
			4584: begin
				if(in == 0) begin
					state<=3905;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=7;
					out<=138;
				end
				if(in == 3) begin
					state<=5894;
					out<=139;
				end
				if(in == 4) begin
					state<=2005;
					out<=140;
				end
			end
			4585: begin
				if(in == 0) begin
					state<=3906;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=8;
					out<=143;
				end
				if(in == 3) begin
					state<=5895;
					out<=144;
				end
				if(in == 4) begin
					state<=2006;
					out<=145;
				end
			end
			4586: begin
				if(in == 0) begin
					state<=3907;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=9;
					out<=148;
				end
				if(in == 3) begin
					state<=5896;
					out<=149;
				end
				if(in == 4) begin
					state<=2007;
					out<=150;
				end
			end
			4587: begin
				if(in == 0) begin
					state<=3908;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=10;
					out<=153;
				end
				if(in == 3) begin
					state<=5897;
					out<=154;
				end
				if(in == 4) begin
					state<=2008;
					out<=155;
				end
			end
			4588: begin
				if(in == 0) begin
					state<=3899;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=1;
					out<=158;
				end
				if(in == 3) begin
					state<=5888;
					out<=159;
				end
				if(in == 4) begin
					state<=1999;
					out<=160;
				end
			end
			4589: begin
				if(in == 0) begin
					state<=4600;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=702;
					out<=163;
				end
				if(in == 3) begin
					state<=6589;
					out<=164;
				end
				if(in == 4) begin
					state<=2700;
					out<=165;
				end
			end
			4590: begin
				if(in == 0) begin
					state<=4601;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=703;
					out<=168;
				end
				if(in == 3) begin
					state<=6590;
					out<=169;
				end
				if(in == 4) begin
					state<=2701;
					out<=170;
				end
			end
			4591: begin
				if(in == 0) begin
					state<=4602;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=704;
					out<=173;
				end
				if(in == 3) begin
					state<=6591;
					out<=174;
				end
				if(in == 4) begin
					state<=2702;
					out<=175;
				end
			end
			4592: begin
				if(in == 0) begin
					state<=4603;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=705;
					out<=178;
				end
				if(in == 3) begin
					state<=6592;
					out<=179;
				end
				if(in == 4) begin
					state<=2703;
					out<=180;
				end
			end
			4593: begin
				if(in == 0) begin
					state<=4604;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=706;
					out<=183;
				end
				if(in == 3) begin
					state<=6593;
					out<=184;
				end
				if(in == 4) begin
					state<=2704;
					out<=185;
				end
			end
			4594: begin
				if(in == 0) begin
					state<=4605;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=707;
					out<=188;
				end
				if(in == 3) begin
					state<=6594;
					out<=189;
				end
				if(in == 4) begin
					state<=2705;
					out<=190;
				end
			end
			4595: begin
				if(in == 0) begin
					state<=4606;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=708;
					out<=193;
				end
				if(in == 3) begin
					state<=6595;
					out<=194;
				end
				if(in == 4) begin
					state<=2706;
					out<=195;
				end
			end
			4596: begin
				if(in == 0) begin
					state<=4607;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=709;
					out<=198;
				end
				if(in == 3) begin
					state<=6596;
					out<=199;
				end
				if(in == 4) begin
					state<=2707;
					out<=200;
				end
			end
			4597: begin
				if(in == 0) begin
					state<=4598;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=700;
					out<=203;
				end
				if(in == 3) begin
					state<=6587;
					out<=204;
				end
				if(in == 4) begin
					state<=2698;
					out<=205;
				end
			end
			4598: begin
				if(in == 0) begin
					state<=4609;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=711;
					out<=208;
				end
				if(in == 3) begin
					state<=6598;
					out<=209;
				end
				if(in == 4) begin
					state<=2709;
					out<=210;
				end
			end
			4599: begin
				if(in == 0) begin
					state<=4610;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=712;
					out<=213;
				end
				if(in == 3) begin
					state<=6599;
					out<=214;
				end
				if(in == 4) begin
					state<=2710;
					out<=215;
				end
			end
			4600: begin
				if(in == 0) begin
					state<=4611;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=713;
					out<=218;
				end
				if(in == 3) begin
					state<=6600;
					out<=219;
				end
				if(in == 4) begin
					state<=2711;
					out<=220;
				end
			end
			4601: begin
				if(in == 0) begin
					state<=4612;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=714;
					out<=223;
				end
				if(in == 3) begin
					state<=6601;
					out<=224;
				end
				if(in == 4) begin
					state<=2712;
					out<=225;
				end
			end
			4602: begin
				if(in == 0) begin
					state<=4613;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=715;
					out<=228;
				end
				if(in == 3) begin
					state<=6602;
					out<=229;
				end
				if(in == 4) begin
					state<=2713;
					out<=230;
				end
			end
			4603: begin
				if(in == 0) begin
					state<=4614;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=716;
					out<=233;
				end
				if(in == 3) begin
					state<=6603;
					out<=234;
				end
				if(in == 4) begin
					state<=2714;
					out<=235;
				end
			end
			4604: begin
				if(in == 0) begin
					state<=4615;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=717;
					out<=238;
				end
				if(in == 3) begin
					state<=6604;
					out<=239;
				end
				if(in == 4) begin
					state<=2715;
					out<=240;
				end
			end
			4605: begin
				if(in == 0) begin
					state<=4616;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=718;
					out<=243;
				end
				if(in == 3) begin
					state<=6605;
					out<=244;
				end
				if(in == 4) begin
					state<=2716;
					out<=245;
				end
			end
			4606: begin
				if(in == 0) begin
					state<=4617;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=719;
					out<=248;
				end
				if(in == 3) begin
					state<=6606;
					out<=249;
				end
				if(in == 4) begin
					state<=2717;
					out<=250;
				end
			end
			4607: begin
				if(in == 0) begin
					state<=4608;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=710;
					out<=253;
				end
				if(in == 3) begin
					state<=6597;
					out<=254;
				end
				if(in == 4) begin
					state<=2708;
					out<=255;
				end
			end
			4608: begin
				if(in == 0) begin
					state<=4619;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=721;
					out<=2;
				end
				if(in == 3) begin
					state<=6608;
					out<=3;
				end
				if(in == 4) begin
					state<=2719;
					out<=4;
				end
			end
			4609: begin
				if(in == 0) begin
					state<=4620;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=722;
					out<=7;
				end
				if(in == 3) begin
					state<=6609;
					out<=8;
				end
				if(in == 4) begin
					state<=2720;
					out<=9;
				end
			end
			4610: begin
				if(in == 0) begin
					state<=4621;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=723;
					out<=12;
				end
				if(in == 3) begin
					state<=6610;
					out<=13;
				end
				if(in == 4) begin
					state<=2721;
					out<=14;
				end
			end
			4611: begin
				if(in == 0) begin
					state<=4622;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=724;
					out<=17;
				end
				if(in == 3) begin
					state<=6611;
					out<=18;
				end
				if(in == 4) begin
					state<=2722;
					out<=19;
				end
			end
			4612: begin
				if(in == 0) begin
					state<=4623;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=725;
					out<=22;
				end
				if(in == 3) begin
					state<=6612;
					out<=23;
				end
				if(in == 4) begin
					state<=2723;
					out<=24;
				end
			end
			4613: begin
				if(in == 0) begin
					state<=4624;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=726;
					out<=27;
				end
				if(in == 3) begin
					state<=6613;
					out<=28;
				end
				if(in == 4) begin
					state<=2724;
					out<=29;
				end
			end
			4614: begin
				if(in == 0) begin
					state<=4625;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=727;
					out<=32;
				end
				if(in == 3) begin
					state<=6614;
					out<=33;
				end
				if(in == 4) begin
					state<=2725;
					out<=34;
				end
			end
			4615: begin
				if(in == 0) begin
					state<=4626;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=728;
					out<=37;
				end
				if(in == 3) begin
					state<=6615;
					out<=38;
				end
				if(in == 4) begin
					state<=2726;
					out<=39;
				end
			end
			4616: begin
				if(in == 0) begin
					state<=4627;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=729;
					out<=42;
				end
				if(in == 3) begin
					state<=6616;
					out<=43;
				end
				if(in == 4) begin
					state<=2727;
					out<=44;
				end
			end
			4617: begin
				if(in == 0) begin
					state<=4618;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=720;
					out<=47;
				end
				if(in == 3) begin
					state<=6607;
					out<=48;
				end
				if(in == 4) begin
					state<=2718;
					out<=49;
				end
			end
			4618: begin
				if(in == 0) begin
					state<=4629;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=731;
					out<=52;
				end
				if(in == 3) begin
					state<=6618;
					out<=53;
				end
				if(in == 4) begin
					state<=2729;
					out<=54;
				end
			end
			4619: begin
				if(in == 0) begin
					state<=4630;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=732;
					out<=57;
				end
				if(in == 3) begin
					state<=6619;
					out<=58;
				end
				if(in == 4) begin
					state<=2730;
					out<=59;
				end
			end
			4620: begin
				if(in == 0) begin
					state<=4631;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=733;
					out<=62;
				end
				if(in == 3) begin
					state<=6620;
					out<=63;
				end
				if(in == 4) begin
					state<=2731;
					out<=64;
				end
			end
			4621: begin
				if(in == 0) begin
					state<=4632;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=734;
					out<=67;
				end
				if(in == 3) begin
					state<=6621;
					out<=68;
				end
				if(in == 4) begin
					state<=2732;
					out<=69;
				end
			end
			4622: begin
				if(in == 0) begin
					state<=4633;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=735;
					out<=72;
				end
				if(in == 3) begin
					state<=6622;
					out<=73;
				end
				if(in == 4) begin
					state<=2733;
					out<=74;
				end
			end
			4623: begin
				if(in == 0) begin
					state<=4634;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=736;
					out<=77;
				end
				if(in == 3) begin
					state<=6623;
					out<=78;
				end
				if(in == 4) begin
					state<=2734;
					out<=79;
				end
			end
			4624: begin
				if(in == 0) begin
					state<=4635;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=737;
					out<=82;
				end
				if(in == 3) begin
					state<=6624;
					out<=83;
				end
				if(in == 4) begin
					state<=2735;
					out<=84;
				end
			end
			4625: begin
				if(in == 0) begin
					state<=4636;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=738;
					out<=87;
				end
				if(in == 3) begin
					state<=6625;
					out<=88;
				end
				if(in == 4) begin
					state<=2736;
					out<=89;
				end
			end
			4626: begin
				if(in == 0) begin
					state<=4637;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=739;
					out<=92;
				end
				if(in == 3) begin
					state<=6626;
					out<=93;
				end
				if(in == 4) begin
					state<=2737;
					out<=94;
				end
			end
			4627: begin
				if(in == 0) begin
					state<=4628;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=730;
					out<=97;
				end
				if(in == 3) begin
					state<=6617;
					out<=98;
				end
				if(in == 4) begin
					state<=2728;
					out<=99;
				end
			end
			4628: begin
				if(in == 0) begin
					state<=4639;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=741;
					out<=102;
				end
				if(in == 3) begin
					state<=6628;
					out<=103;
				end
				if(in == 4) begin
					state<=2739;
					out<=104;
				end
			end
			4629: begin
				if(in == 0) begin
					state<=4640;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=742;
					out<=107;
				end
				if(in == 3) begin
					state<=6629;
					out<=108;
				end
				if(in == 4) begin
					state<=2740;
					out<=109;
				end
			end
			4630: begin
				if(in == 0) begin
					state<=4641;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=743;
					out<=112;
				end
				if(in == 3) begin
					state<=6630;
					out<=113;
				end
				if(in == 4) begin
					state<=2741;
					out<=114;
				end
			end
			4631: begin
				if(in == 0) begin
					state<=4642;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=744;
					out<=117;
				end
				if(in == 3) begin
					state<=6631;
					out<=118;
				end
				if(in == 4) begin
					state<=2742;
					out<=119;
				end
			end
			4632: begin
				if(in == 0) begin
					state<=4643;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=745;
					out<=122;
				end
				if(in == 3) begin
					state<=6632;
					out<=123;
				end
				if(in == 4) begin
					state<=2743;
					out<=124;
				end
			end
			4633: begin
				if(in == 0) begin
					state<=4644;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=746;
					out<=127;
				end
				if(in == 3) begin
					state<=6633;
					out<=128;
				end
				if(in == 4) begin
					state<=2744;
					out<=129;
				end
			end
			4634: begin
				if(in == 0) begin
					state<=4645;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=747;
					out<=132;
				end
				if(in == 3) begin
					state<=6634;
					out<=133;
				end
				if(in == 4) begin
					state<=2745;
					out<=134;
				end
			end
			4635: begin
				if(in == 0) begin
					state<=4646;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=748;
					out<=137;
				end
				if(in == 3) begin
					state<=6635;
					out<=138;
				end
				if(in == 4) begin
					state<=2746;
					out<=139;
				end
			end
			4636: begin
				if(in == 0) begin
					state<=4647;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=749;
					out<=142;
				end
				if(in == 3) begin
					state<=6636;
					out<=143;
				end
				if(in == 4) begin
					state<=2747;
					out<=144;
				end
			end
			4637: begin
				if(in == 0) begin
					state<=4638;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=740;
					out<=147;
				end
				if(in == 3) begin
					state<=6627;
					out<=148;
				end
				if(in == 4) begin
					state<=2738;
					out<=149;
				end
			end
			4638: begin
				if(in == 0) begin
					state<=4649;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=751;
					out<=152;
				end
				if(in == 3) begin
					state<=6638;
					out<=153;
				end
				if(in == 4) begin
					state<=2749;
					out<=154;
				end
			end
			4639: begin
				if(in == 0) begin
					state<=4650;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=752;
					out<=157;
				end
				if(in == 3) begin
					state<=6639;
					out<=158;
				end
				if(in == 4) begin
					state<=2750;
					out<=159;
				end
			end
			4640: begin
				if(in == 0) begin
					state<=4651;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=753;
					out<=162;
				end
				if(in == 3) begin
					state<=6640;
					out<=163;
				end
				if(in == 4) begin
					state<=2751;
					out<=164;
				end
			end
			4641: begin
				if(in == 0) begin
					state<=4652;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=754;
					out<=167;
				end
				if(in == 3) begin
					state<=6641;
					out<=168;
				end
				if(in == 4) begin
					state<=2752;
					out<=169;
				end
			end
			4642: begin
				if(in == 0) begin
					state<=4653;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=755;
					out<=172;
				end
				if(in == 3) begin
					state<=6642;
					out<=173;
				end
				if(in == 4) begin
					state<=2753;
					out<=174;
				end
			end
			4643: begin
				if(in == 0) begin
					state<=4654;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=756;
					out<=177;
				end
				if(in == 3) begin
					state<=6643;
					out<=178;
				end
				if(in == 4) begin
					state<=2754;
					out<=179;
				end
			end
			4644: begin
				if(in == 0) begin
					state<=4655;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=757;
					out<=182;
				end
				if(in == 3) begin
					state<=6644;
					out<=183;
				end
				if(in == 4) begin
					state<=2755;
					out<=184;
				end
			end
			4645: begin
				if(in == 0) begin
					state<=4656;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=758;
					out<=187;
				end
				if(in == 3) begin
					state<=6645;
					out<=188;
				end
				if(in == 4) begin
					state<=2756;
					out<=189;
				end
			end
			4646: begin
				if(in == 0) begin
					state<=4657;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=759;
					out<=192;
				end
				if(in == 3) begin
					state<=6646;
					out<=193;
				end
				if(in == 4) begin
					state<=2757;
					out<=194;
				end
			end
			4647: begin
				if(in == 0) begin
					state<=4648;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=750;
					out<=197;
				end
				if(in == 3) begin
					state<=6637;
					out<=198;
				end
				if(in == 4) begin
					state<=2748;
					out<=199;
				end
			end
			4648: begin
				if(in == 0) begin
					state<=4659;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=761;
					out<=202;
				end
				if(in == 3) begin
					state<=6648;
					out<=203;
				end
				if(in == 4) begin
					state<=2759;
					out<=204;
				end
			end
			4649: begin
				if(in == 0) begin
					state<=4660;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=762;
					out<=207;
				end
				if(in == 3) begin
					state<=6649;
					out<=208;
				end
				if(in == 4) begin
					state<=2760;
					out<=209;
				end
			end
			4650: begin
				if(in == 0) begin
					state<=4661;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=763;
					out<=212;
				end
				if(in == 3) begin
					state<=6650;
					out<=213;
				end
				if(in == 4) begin
					state<=2761;
					out<=214;
				end
			end
			4651: begin
				if(in == 0) begin
					state<=4662;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=764;
					out<=217;
				end
				if(in == 3) begin
					state<=6651;
					out<=218;
				end
				if(in == 4) begin
					state<=2762;
					out<=219;
				end
			end
			4652: begin
				if(in == 0) begin
					state<=4663;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=765;
					out<=222;
				end
				if(in == 3) begin
					state<=6652;
					out<=223;
				end
				if(in == 4) begin
					state<=2763;
					out<=224;
				end
			end
			4653: begin
				if(in == 0) begin
					state<=4664;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=766;
					out<=227;
				end
				if(in == 3) begin
					state<=6653;
					out<=228;
				end
				if(in == 4) begin
					state<=2764;
					out<=229;
				end
			end
			4654: begin
				if(in == 0) begin
					state<=4665;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=767;
					out<=232;
				end
				if(in == 3) begin
					state<=6654;
					out<=233;
				end
				if(in == 4) begin
					state<=2765;
					out<=234;
				end
			end
			4655: begin
				if(in == 0) begin
					state<=4666;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=768;
					out<=237;
				end
				if(in == 3) begin
					state<=6655;
					out<=238;
				end
				if(in == 4) begin
					state<=2766;
					out<=239;
				end
			end
			4656: begin
				if(in == 0) begin
					state<=4667;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=769;
					out<=242;
				end
				if(in == 3) begin
					state<=6656;
					out<=243;
				end
				if(in == 4) begin
					state<=2767;
					out<=244;
				end
			end
			4657: begin
				if(in == 0) begin
					state<=4658;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=760;
					out<=247;
				end
				if(in == 3) begin
					state<=6647;
					out<=248;
				end
				if(in == 4) begin
					state<=2758;
					out<=249;
				end
			end
			4658: begin
				if(in == 0) begin
					state<=4669;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=771;
					out<=252;
				end
				if(in == 3) begin
					state<=6658;
					out<=253;
				end
				if(in == 4) begin
					state<=2769;
					out<=254;
				end
			end
			4659: begin
				if(in == 0) begin
					state<=4670;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=772;
					out<=1;
				end
				if(in == 3) begin
					state<=6659;
					out<=2;
				end
				if(in == 4) begin
					state<=2770;
					out<=3;
				end
			end
			4660: begin
				if(in == 0) begin
					state<=4671;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=773;
					out<=6;
				end
				if(in == 3) begin
					state<=6660;
					out<=7;
				end
				if(in == 4) begin
					state<=2771;
					out<=8;
				end
			end
			4661: begin
				if(in == 0) begin
					state<=4672;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=774;
					out<=11;
				end
				if(in == 3) begin
					state<=6661;
					out<=12;
				end
				if(in == 4) begin
					state<=2772;
					out<=13;
				end
			end
			4662: begin
				if(in == 0) begin
					state<=4673;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=775;
					out<=16;
				end
				if(in == 3) begin
					state<=6662;
					out<=17;
				end
				if(in == 4) begin
					state<=2773;
					out<=18;
				end
			end
			4663: begin
				if(in == 0) begin
					state<=4674;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=776;
					out<=21;
				end
				if(in == 3) begin
					state<=6663;
					out<=22;
				end
				if(in == 4) begin
					state<=2774;
					out<=23;
				end
			end
			4664: begin
				if(in == 0) begin
					state<=4675;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=777;
					out<=26;
				end
				if(in == 3) begin
					state<=6664;
					out<=27;
				end
				if(in == 4) begin
					state<=2775;
					out<=28;
				end
			end
			4665: begin
				if(in == 0) begin
					state<=4676;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=778;
					out<=31;
				end
				if(in == 3) begin
					state<=6665;
					out<=32;
				end
				if(in == 4) begin
					state<=2776;
					out<=33;
				end
			end
			4666: begin
				if(in == 0) begin
					state<=4677;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=779;
					out<=36;
				end
				if(in == 3) begin
					state<=6666;
					out<=37;
				end
				if(in == 4) begin
					state<=2777;
					out<=38;
				end
			end
			4667: begin
				if(in == 0) begin
					state<=4668;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=770;
					out<=41;
				end
				if(in == 3) begin
					state<=6657;
					out<=42;
				end
				if(in == 4) begin
					state<=2768;
					out<=43;
				end
			end
			4668: begin
				if(in == 0) begin
					state<=4679;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=781;
					out<=46;
				end
				if(in == 3) begin
					state<=6668;
					out<=47;
				end
				if(in == 4) begin
					state<=2779;
					out<=48;
				end
			end
			4669: begin
				if(in == 0) begin
					state<=4680;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=782;
					out<=51;
				end
				if(in == 3) begin
					state<=6669;
					out<=52;
				end
				if(in == 4) begin
					state<=2780;
					out<=53;
				end
			end
			4670: begin
				if(in == 0) begin
					state<=4681;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=783;
					out<=56;
				end
				if(in == 3) begin
					state<=6670;
					out<=57;
				end
				if(in == 4) begin
					state<=2781;
					out<=58;
				end
			end
			4671: begin
				if(in == 0) begin
					state<=4682;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=784;
					out<=61;
				end
				if(in == 3) begin
					state<=6671;
					out<=62;
				end
				if(in == 4) begin
					state<=2782;
					out<=63;
				end
			end
			4672: begin
				if(in == 0) begin
					state<=4683;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=785;
					out<=66;
				end
				if(in == 3) begin
					state<=6672;
					out<=67;
				end
				if(in == 4) begin
					state<=2783;
					out<=68;
				end
			end
			4673: begin
				if(in == 0) begin
					state<=4684;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=786;
					out<=71;
				end
				if(in == 3) begin
					state<=6673;
					out<=72;
				end
				if(in == 4) begin
					state<=2784;
					out<=73;
				end
			end
			4674: begin
				if(in == 0) begin
					state<=4685;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=787;
					out<=76;
				end
				if(in == 3) begin
					state<=6674;
					out<=77;
				end
				if(in == 4) begin
					state<=2785;
					out<=78;
				end
			end
			4675: begin
				if(in == 0) begin
					state<=4686;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=788;
					out<=81;
				end
				if(in == 3) begin
					state<=6675;
					out<=82;
				end
				if(in == 4) begin
					state<=2786;
					out<=83;
				end
			end
			4676: begin
				if(in == 0) begin
					state<=4687;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=789;
					out<=86;
				end
				if(in == 3) begin
					state<=6676;
					out<=87;
				end
				if(in == 4) begin
					state<=2787;
					out<=88;
				end
			end
			4677: begin
				if(in == 0) begin
					state<=4678;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=780;
					out<=91;
				end
				if(in == 3) begin
					state<=6667;
					out<=92;
				end
				if(in == 4) begin
					state<=2778;
					out<=93;
				end
			end
			4678: begin
				if(in == 0) begin
					state<=4689;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=791;
					out<=96;
				end
				if(in == 3) begin
					state<=6678;
					out<=97;
				end
				if(in == 4) begin
					state<=2789;
					out<=98;
				end
			end
			4679: begin
				if(in == 0) begin
					state<=4690;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=792;
					out<=101;
				end
				if(in == 3) begin
					state<=6679;
					out<=102;
				end
				if(in == 4) begin
					state<=2790;
					out<=103;
				end
			end
			4680: begin
				if(in == 0) begin
					state<=4691;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=793;
					out<=106;
				end
				if(in == 3) begin
					state<=6680;
					out<=107;
				end
				if(in == 4) begin
					state<=2791;
					out<=108;
				end
			end
			4681: begin
				if(in == 0) begin
					state<=4692;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=794;
					out<=111;
				end
				if(in == 3) begin
					state<=6681;
					out<=112;
				end
				if(in == 4) begin
					state<=2792;
					out<=113;
				end
			end
			4682: begin
				if(in == 0) begin
					state<=4693;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=795;
					out<=116;
				end
				if(in == 3) begin
					state<=6682;
					out<=117;
				end
				if(in == 4) begin
					state<=2793;
					out<=118;
				end
			end
			4683: begin
				if(in == 0) begin
					state<=4694;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=796;
					out<=121;
				end
				if(in == 3) begin
					state<=6683;
					out<=122;
				end
				if(in == 4) begin
					state<=2794;
					out<=123;
				end
			end
			4684: begin
				if(in == 0) begin
					state<=4695;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=797;
					out<=126;
				end
				if(in == 3) begin
					state<=6684;
					out<=127;
				end
				if(in == 4) begin
					state<=2795;
					out<=128;
				end
			end
			4685: begin
				if(in == 0) begin
					state<=4696;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=798;
					out<=131;
				end
				if(in == 3) begin
					state<=6685;
					out<=132;
				end
				if(in == 4) begin
					state<=2796;
					out<=133;
				end
			end
			4686: begin
				if(in == 0) begin
					state<=4697;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=799;
					out<=136;
				end
				if(in == 3) begin
					state<=6686;
					out<=137;
				end
				if(in == 4) begin
					state<=2797;
					out<=138;
				end
			end
			4687: begin
				if(in == 0) begin
					state<=4688;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=790;
					out<=141;
				end
				if(in == 3) begin
					state<=6677;
					out<=142;
				end
				if(in == 4) begin
					state<=2788;
					out<=143;
				end
			end
			4688: begin
				if(in == 0) begin
					state<=4709;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=811;
					out<=146;
				end
				if(in == 3) begin
					state<=6698;
					out<=147;
				end
				if(in == 4) begin
					state<=2809;
					out<=148;
				end
			end
			4689: begin
				if(in == 0) begin
					state<=4710;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=812;
					out<=151;
				end
				if(in == 3) begin
					state<=6699;
					out<=152;
				end
				if(in == 4) begin
					state<=2810;
					out<=153;
				end
			end
			4690: begin
				if(in == 0) begin
					state<=4711;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=813;
					out<=156;
				end
				if(in == 3) begin
					state<=6700;
					out<=157;
				end
				if(in == 4) begin
					state<=2811;
					out<=158;
				end
			end
			4691: begin
				if(in == 0) begin
					state<=4712;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=814;
					out<=161;
				end
				if(in == 3) begin
					state<=6701;
					out<=162;
				end
				if(in == 4) begin
					state<=2812;
					out<=163;
				end
			end
			4692: begin
				if(in == 0) begin
					state<=4713;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=815;
					out<=166;
				end
				if(in == 3) begin
					state<=6702;
					out<=167;
				end
				if(in == 4) begin
					state<=2813;
					out<=168;
				end
			end
			4693: begin
				if(in == 0) begin
					state<=4714;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=816;
					out<=171;
				end
				if(in == 3) begin
					state<=6703;
					out<=172;
				end
				if(in == 4) begin
					state<=2814;
					out<=173;
				end
			end
			4694: begin
				if(in == 0) begin
					state<=4715;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=817;
					out<=176;
				end
				if(in == 3) begin
					state<=6704;
					out<=177;
				end
				if(in == 4) begin
					state<=2815;
					out<=178;
				end
			end
			4695: begin
				if(in == 0) begin
					state<=4716;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=818;
					out<=181;
				end
				if(in == 3) begin
					state<=6705;
					out<=182;
				end
				if(in == 4) begin
					state<=2816;
					out<=183;
				end
			end
			4696: begin
				if(in == 0) begin
					state<=4717;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=819;
					out<=186;
				end
				if(in == 3) begin
					state<=6706;
					out<=187;
				end
				if(in == 4) begin
					state<=2817;
					out<=188;
				end
			end
			4697: begin
				if(in == 0) begin
					state<=4708;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=810;
					out<=191;
				end
				if(in == 3) begin
					state<=6697;
					out<=192;
				end
				if(in == 4) begin
					state<=2808;
					out<=193;
				end
			end
			4698: begin
				if(in == 0) begin
					state<=5498;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=1609;
					out<=196;
				end
				if(in == 3) begin
					state<=7399;
					out<=197;
				end
				if(in == 4) begin
					state<=3510;
					out<=198;
				end
			end
			4699: begin
				if(in == 0) begin
					state<=5499;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=1610;
					out<=201;
				end
				if(in == 3) begin
					state<=7400;
					out<=202;
				end
				if(in == 4) begin
					state<=3511;
					out<=203;
				end
			end
			4700: begin
				if(in == 0) begin
					state<=5500;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=1611;
					out<=206;
				end
				if(in == 3) begin
					state<=7401;
					out<=207;
				end
				if(in == 4) begin
					state<=3512;
					out<=208;
				end
			end
			4701: begin
				if(in == 0) begin
					state<=5501;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=1612;
					out<=211;
				end
				if(in == 3) begin
					state<=7402;
					out<=212;
				end
				if(in == 4) begin
					state<=3513;
					out<=213;
				end
			end
			4702: begin
				if(in == 0) begin
					state<=5502;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=1613;
					out<=216;
				end
				if(in == 3) begin
					state<=7403;
					out<=217;
				end
				if(in == 4) begin
					state<=3514;
					out<=218;
				end
			end
			4703: begin
				if(in == 0) begin
					state<=5503;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=1614;
					out<=221;
				end
				if(in == 3) begin
					state<=7404;
					out<=222;
				end
				if(in == 4) begin
					state<=3515;
					out<=223;
				end
			end
			4704: begin
				if(in == 0) begin
					state<=5504;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=1615;
					out<=226;
				end
				if(in == 3) begin
					state<=7405;
					out<=227;
				end
				if(in == 4) begin
					state<=3516;
					out<=228;
				end
			end
			4705: begin
				if(in == 0) begin
					state<=5505;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=1616;
					out<=231;
				end
				if(in == 3) begin
					state<=7406;
					out<=232;
				end
				if(in == 4) begin
					state<=3517;
					out<=233;
				end
			end
			4706: begin
				if(in == 0) begin
					state<=5506;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=1617;
					out<=236;
				end
				if(in == 3) begin
					state<=7407;
					out<=237;
				end
				if(in == 4) begin
					state<=3518;
					out<=238;
				end
			end
			4707: begin
				if(in == 0) begin
					state<=5497;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=1608;
					out<=241;
				end
				if(in == 3) begin
					state<=7398;
					out<=242;
				end
				if(in == 4) begin
					state<=3509;
					out<=243;
				end
			end
			4708: begin
				if(in == 0) begin
					state<=4719;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=821;
					out<=246;
				end
				if(in == 3) begin
					state<=6708;
					out<=247;
				end
				if(in == 4) begin
					state<=2819;
					out<=248;
				end
			end
			4709: begin
				if(in == 0) begin
					state<=4720;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=822;
					out<=251;
				end
				if(in == 3) begin
					state<=6709;
					out<=252;
				end
				if(in == 4) begin
					state<=2820;
					out<=253;
				end
			end
			4710: begin
				if(in == 0) begin
					state<=4721;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=823;
					out<=0;
				end
				if(in == 3) begin
					state<=6710;
					out<=1;
				end
				if(in == 4) begin
					state<=2821;
					out<=2;
				end
			end
			4711: begin
				if(in == 0) begin
					state<=4722;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=824;
					out<=5;
				end
				if(in == 3) begin
					state<=6711;
					out<=6;
				end
				if(in == 4) begin
					state<=2822;
					out<=7;
				end
			end
			4712: begin
				if(in == 0) begin
					state<=4723;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=825;
					out<=10;
				end
				if(in == 3) begin
					state<=6712;
					out<=11;
				end
				if(in == 4) begin
					state<=2823;
					out<=12;
				end
			end
			4713: begin
				if(in == 0) begin
					state<=4724;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=826;
					out<=15;
				end
				if(in == 3) begin
					state<=6713;
					out<=16;
				end
				if(in == 4) begin
					state<=2824;
					out<=17;
				end
			end
			4714: begin
				if(in == 0) begin
					state<=4725;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=827;
					out<=20;
				end
				if(in == 3) begin
					state<=6714;
					out<=21;
				end
				if(in == 4) begin
					state<=2825;
					out<=22;
				end
			end
			4715: begin
				if(in == 0) begin
					state<=4726;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=828;
					out<=25;
				end
				if(in == 3) begin
					state<=6715;
					out<=26;
				end
				if(in == 4) begin
					state<=2826;
					out<=27;
				end
			end
			4716: begin
				if(in == 0) begin
					state<=4727;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=829;
					out<=30;
				end
				if(in == 3) begin
					state<=6716;
					out<=31;
				end
				if(in == 4) begin
					state<=2827;
					out<=32;
				end
			end
			4717: begin
				if(in == 0) begin
					state<=4718;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=820;
					out<=35;
				end
				if(in == 3) begin
					state<=6707;
					out<=36;
				end
				if(in == 4) begin
					state<=2818;
					out<=37;
				end
			end
			4718: begin
				if(in == 0) begin
					state<=4729;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=831;
					out<=40;
				end
				if(in == 3) begin
					state<=6718;
					out<=41;
				end
				if(in == 4) begin
					state<=2829;
					out<=42;
				end
			end
			4719: begin
				if(in == 0) begin
					state<=4730;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=832;
					out<=45;
				end
				if(in == 3) begin
					state<=6719;
					out<=46;
				end
				if(in == 4) begin
					state<=2830;
					out<=47;
				end
			end
			4720: begin
				if(in == 0) begin
					state<=4731;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=833;
					out<=50;
				end
				if(in == 3) begin
					state<=6720;
					out<=51;
				end
				if(in == 4) begin
					state<=2831;
					out<=52;
				end
			end
			4721: begin
				if(in == 0) begin
					state<=4732;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=834;
					out<=55;
				end
				if(in == 3) begin
					state<=6721;
					out<=56;
				end
				if(in == 4) begin
					state<=2832;
					out<=57;
				end
			end
			4722: begin
				if(in == 0) begin
					state<=4733;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=835;
					out<=60;
				end
				if(in == 3) begin
					state<=6722;
					out<=61;
				end
				if(in == 4) begin
					state<=2833;
					out<=62;
				end
			end
			4723: begin
				if(in == 0) begin
					state<=4734;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=836;
					out<=65;
				end
				if(in == 3) begin
					state<=6723;
					out<=66;
				end
				if(in == 4) begin
					state<=2834;
					out<=67;
				end
			end
			4724: begin
				if(in == 0) begin
					state<=4735;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=837;
					out<=70;
				end
				if(in == 3) begin
					state<=6724;
					out<=71;
				end
				if(in == 4) begin
					state<=2835;
					out<=72;
				end
			end
			4725: begin
				if(in == 0) begin
					state<=4736;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=838;
					out<=75;
				end
				if(in == 3) begin
					state<=6725;
					out<=76;
				end
				if(in == 4) begin
					state<=2836;
					out<=77;
				end
			end
			4726: begin
				if(in == 0) begin
					state<=4737;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=839;
					out<=80;
				end
				if(in == 3) begin
					state<=6726;
					out<=81;
				end
				if(in == 4) begin
					state<=2837;
					out<=82;
				end
			end
			4727: begin
				if(in == 0) begin
					state<=4728;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=830;
					out<=85;
				end
				if(in == 3) begin
					state<=6717;
					out<=86;
				end
				if(in == 4) begin
					state<=2828;
					out<=87;
				end
			end
			4728: begin
				if(in == 0) begin
					state<=4739;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=841;
					out<=90;
				end
				if(in == 3) begin
					state<=6728;
					out<=91;
				end
				if(in == 4) begin
					state<=2839;
					out<=92;
				end
			end
			4729: begin
				if(in == 0) begin
					state<=4740;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=842;
					out<=95;
				end
				if(in == 3) begin
					state<=6729;
					out<=96;
				end
				if(in == 4) begin
					state<=2840;
					out<=97;
				end
			end
			4730: begin
				if(in == 0) begin
					state<=4741;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=843;
					out<=100;
				end
				if(in == 3) begin
					state<=6730;
					out<=101;
				end
				if(in == 4) begin
					state<=2841;
					out<=102;
				end
			end
			4731: begin
				if(in == 0) begin
					state<=4742;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=844;
					out<=105;
				end
				if(in == 3) begin
					state<=6731;
					out<=106;
				end
				if(in == 4) begin
					state<=2842;
					out<=107;
				end
			end
			4732: begin
				if(in == 0) begin
					state<=4743;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=845;
					out<=110;
				end
				if(in == 3) begin
					state<=6732;
					out<=111;
				end
				if(in == 4) begin
					state<=2843;
					out<=112;
				end
			end
			4733: begin
				if(in == 0) begin
					state<=4744;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=846;
					out<=115;
				end
				if(in == 3) begin
					state<=6733;
					out<=116;
				end
				if(in == 4) begin
					state<=2844;
					out<=117;
				end
			end
			4734: begin
				if(in == 0) begin
					state<=4745;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=847;
					out<=120;
				end
				if(in == 3) begin
					state<=6734;
					out<=121;
				end
				if(in == 4) begin
					state<=2845;
					out<=122;
				end
			end
			4735: begin
				if(in == 0) begin
					state<=4746;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=848;
					out<=125;
				end
				if(in == 3) begin
					state<=6735;
					out<=126;
				end
				if(in == 4) begin
					state<=2846;
					out<=127;
				end
			end
			4736: begin
				if(in == 0) begin
					state<=4747;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=849;
					out<=130;
				end
				if(in == 3) begin
					state<=6736;
					out<=131;
				end
				if(in == 4) begin
					state<=2847;
					out<=132;
				end
			end
			4737: begin
				if(in == 0) begin
					state<=4738;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=840;
					out<=135;
				end
				if(in == 3) begin
					state<=6727;
					out<=136;
				end
				if(in == 4) begin
					state<=2838;
					out<=137;
				end
			end
			4738: begin
				if(in == 0) begin
					state<=4749;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=851;
					out<=140;
				end
				if(in == 3) begin
					state<=6738;
					out<=141;
				end
				if(in == 4) begin
					state<=2849;
					out<=142;
				end
			end
			4739: begin
				if(in == 0) begin
					state<=4750;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=852;
					out<=145;
				end
				if(in == 3) begin
					state<=6739;
					out<=146;
				end
				if(in == 4) begin
					state<=2850;
					out<=147;
				end
			end
			4740: begin
				if(in == 0) begin
					state<=4751;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=853;
					out<=150;
				end
				if(in == 3) begin
					state<=6740;
					out<=151;
				end
				if(in == 4) begin
					state<=2851;
					out<=152;
				end
			end
			4741: begin
				if(in == 0) begin
					state<=4752;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=854;
					out<=155;
				end
				if(in == 3) begin
					state<=6741;
					out<=156;
				end
				if(in == 4) begin
					state<=2852;
					out<=157;
				end
			end
			4742: begin
				if(in == 0) begin
					state<=4753;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=855;
					out<=160;
				end
				if(in == 3) begin
					state<=6742;
					out<=161;
				end
				if(in == 4) begin
					state<=2853;
					out<=162;
				end
			end
			4743: begin
				if(in == 0) begin
					state<=4754;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=856;
					out<=165;
				end
				if(in == 3) begin
					state<=6743;
					out<=166;
				end
				if(in == 4) begin
					state<=2854;
					out<=167;
				end
			end
			4744: begin
				if(in == 0) begin
					state<=4755;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=857;
					out<=170;
				end
				if(in == 3) begin
					state<=6744;
					out<=171;
				end
				if(in == 4) begin
					state<=2855;
					out<=172;
				end
			end
			4745: begin
				if(in == 0) begin
					state<=4756;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=858;
					out<=175;
				end
				if(in == 3) begin
					state<=6745;
					out<=176;
				end
				if(in == 4) begin
					state<=2856;
					out<=177;
				end
			end
			4746: begin
				if(in == 0) begin
					state<=4757;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=859;
					out<=180;
				end
				if(in == 3) begin
					state<=6746;
					out<=181;
				end
				if(in == 4) begin
					state<=2857;
					out<=182;
				end
			end
			4747: begin
				if(in == 0) begin
					state<=4748;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=850;
					out<=185;
				end
				if(in == 3) begin
					state<=6737;
					out<=186;
				end
				if(in == 4) begin
					state<=2848;
					out<=187;
				end
			end
			4748: begin
				if(in == 0) begin
					state<=4759;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=861;
					out<=190;
				end
				if(in == 3) begin
					state<=6748;
					out<=191;
				end
				if(in == 4) begin
					state<=2859;
					out<=192;
				end
			end
			4749: begin
				if(in == 0) begin
					state<=4760;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=862;
					out<=195;
				end
				if(in == 3) begin
					state<=6749;
					out<=196;
				end
				if(in == 4) begin
					state<=2860;
					out<=197;
				end
			end
			4750: begin
				if(in == 0) begin
					state<=4761;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=863;
					out<=200;
				end
				if(in == 3) begin
					state<=6750;
					out<=201;
				end
				if(in == 4) begin
					state<=2861;
					out<=202;
				end
			end
			4751: begin
				if(in == 0) begin
					state<=4762;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=864;
					out<=205;
				end
				if(in == 3) begin
					state<=6751;
					out<=206;
				end
				if(in == 4) begin
					state<=2862;
					out<=207;
				end
			end
			4752: begin
				if(in == 0) begin
					state<=4763;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=865;
					out<=210;
				end
				if(in == 3) begin
					state<=6752;
					out<=211;
				end
				if(in == 4) begin
					state<=2863;
					out<=212;
				end
			end
			4753: begin
				if(in == 0) begin
					state<=4764;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=866;
					out<=215;
				end
				if(in == 3) begin
					state<=6753;
					out<=216;
				end
				if(in == 4) begin
					state<=2864;
					out<=217;
				end
			end
			4754: begin
				if(in == 0) begin
					state<=4765;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=867;
					out<=220;
				end
				if(in == 3) begin
					state<=6754;
					out<=221;
				end
				if(in == 4) begin
					state<=2865;
					out<=222;
				end
			end
			4755: begin
				if(in == 0) begin
					state<=4766;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=868;
					out<=225;
				end
				if(in == 3) begin
					state<=6755;
					out<=226;
				end
				if(in == 4) begin
					state<=2866;
					out<=227;
				end
			end
			4756: begin
				if(in == 0) begin
					state<=4767;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=869;
					out<=230;
				end
				if(in == 3) begin
					state<=6756;
					out<=231;
				end
				if(in == 4) begin
					state<=2867;
					out<=232;
				end
			end
			4757: begin
				if(in == 0) begin
					state<=4758;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=860;
					out<=235;
				end
				if(in == 3) begin
					state<=6747;
					out<=236;
				end
				if(in == 4) begin
					state<=2858;
					out<=237;
				end
			end
			4758: begin
				if(in == 0) begin
					state<=4769;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=871;
					out<=240;
				end
				if(in == 3) begin
					state<=6758;
					out<=241;
				end
				if(in == 4) begin
					state<=2869;
					out<=242;
				end
			end
			4759: begin
				if(in == 0) begin
					state<=4770;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=872;
					out<=245;
				end
				if(in == 3) begin
					state<=6759;
					out<=246;
				end
				if(in == 4) begin
					state<=2870;
					out<=247;
				end
			end
			4760: begin
				if(in == 0) begin
					state<=4771;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=873;
					out<=250;
				end
				if(in == 3) begin
					state<=6760;
					out<=251;
				end
				if(in == 4) begin
					state<=2871;
					out<=252;
				end
			end
			4761: begin
				if(in == 0) begin
					state<=4772;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=874;
					out<=255;
				end
				if(in == 3) begin
					state<=6761;
					out<=0;
				end
				if(in == 4) begin
					state<=2872;
					out<=1;
				end
			end
			4762: begin
				if(in == 0) begin
					state<=4773;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=875;
					out<=4;
				end
				if(in == 3) begin
					state<=6762;
					out<=5;
				end
				if(in == 4) begin
					state<=2873;
					out<=6;
				end
			end
			4763: begin
				if(in == 0) begin
					state<=4774;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=876;
					out<=9;
				end
				if(in == 3) begin
					state<=6763;
					out<=10;
				end
				if(in == 4) begin
					state<=2874;
					out<=11;
				end
			end
			4764: begin
				if(in == 0) begin
					state<=4775;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=877;
					out<=14;
				end
				if(in == 3) begin
					state<=6764;
					out<=15;
				end
				if(in == 4) begin
					state<=2875;
					out<=16;
				end
			end
			4765: begin
				if(in == 0) begin
					state<=4776;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=878;
					out<=19;
				end
				if(in == 3) begin
					state<=6765;
					out<=20;
				end
				if(in == 4) begin
					state<=2876;
					out<=21;
				end
			end
			4766: begin
				if(in == 0) begin
					state<=4777;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=879;
					out<=24;
				end
				if(in == 3) begin
					state<=6766;
					out<=25;
				end
				if(in == 4) begin
					state<=2877;
					out<=26;
				end
			end
			4767: begin
				if(in == 0) begin
					state<=4768;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=870;
					out<=29;
				end
				if(in == 3) begin
					state<=6757;
					out<=30;
				end
				if(in == 4) begin
					state<=2868;
					out<=31;
				end
			end
			4768: begin
				if(in == 0) begin
					state<=4779;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=881;
					out<=34;
				end
				if(in == 3) begin
					state<=6768;
					out<=35;
				end
				if(in == 4) begin
					state<=2879;
					out<=36;
				end
			end
			4769: begin
				if(in == 0) begin
					state<=4780;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=882;
					out<=39;
				end
				if(in == 3) begin
					state<=6769;
					out<=40;
				end
				if(in == 4) begin
					state<=2880;
					out<=41;
				end
			end
			4770: begin
				if(in == 0) begin
					state<=4781;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=883;
					out<=44;
				end
				if(in == 3) begin
					state<=6770;
					out<=45;
				end
				if(in == 4) begin
					state<=2881;
					out<=46;
				end
			end
			4771: begin
				if(in == 0) begin
					state<=4782;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=884;
					out<=49;
				end
				if(in == 3) begin
					state<=6771;
					out<=50;
				end
				if(in == 4) begin
					state<=2882;
					out<=51;
				end
			end
			4772: begin
				if(in == 0) begin
					state<=4783;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=885;
					out<=54;
				end
				if(in == 3) begin
					state<=6772;
					out<=55;
				end
				if(in == 4) begin
					state<=2883;
					out<=56;
				end
			end
			4773: begin
				if(in == 0) begin
					state<=4784;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=886;
					out<=59;
				end
				if(in == 3) begin
					state<=6773;
					out<=60;
				end
				if(in == 4) begin
					state<=2884;
					out<=61;
				end
			end
			4774: begin
				if(in == 0) begin
					state<=4785;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=887;
					out<=64;
				end
				if(in == 3) begin
					state<=6774;
					out<=65;
				end
				if(in == 4) begin
					state<=2885;
					out<=66;
				end
			end
			4775: begin
				if(in == 0) begin
					state<=4786;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=888;
					out<=69;
				end
				if(in == 3) begin
					state<=6775;
					out<=70;
				end
				if(in == 4) begin
					state<=2886;
					out<=71;
				end
			end
			4776: begin
				if(in == 0) begin
					state<=4787;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=889;
					out<=74;
				end
				if(in == 3) begin
					state<=6776;
					out<=75;
				end
				if(in == 4) begin
					state<=2887;
					out<=76;
				end
			end
			4777: begin
				if(in == 0) begin
					state<=4778;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=880;
					out<=79;
				end
				if(in == 3) begin
					state<=6767;
					out<=80;
				end
				if(in == 4) begin
					state<=2878;
					out<=81;
				end
			end
			4778: begin
				if(in == 0) begin
					state<=4789;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=891;
					out<=84;
				end
				if(in == 3) begin
					state<=6778;
					out<=85;
				end
				if(in == 4) begin
					state<=2889;
					out<=86;
				end
			end
			4779: begin
				if(in == 0) begin
					state<=4790;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=892;
					out<=89;
				end
				if(in == 3) begin
					state<=6779;
					out<=90;
				end
				if(in == 4) begin
					state<=2890;
					out<=91;
				end
			end
			4780: begin
				if(in == 0) begin
					state<=4791;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=893;
					out<=94;
				end
				if(in == 3) begin
					state<=6780;
					out<=95;
				end
				if(in == 4) begin
					state<=2891;
					out<=96;
				end
			end
			4781: begin
				if(in == 0) begin
					state<=4792;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=894;
					out<=99;
				end
				if(in == 3) begin
					state<=6781;
					out<=100;
				end
				if(in == 4) begin
					state<=2892;
					out<=101;
				end
			end
			4782: begin
				if(in == 0) begin
					state<=4793;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=895;
					out<=104;
				end
				if(in == 3) begin
					state<=6782;
					out<=105;
				end
				if(in == 4) begin
					state<=2893;
					out<=106;
				end
			end
			4783: begin
				if(in == 0) begin
					state<=4794;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=896;
					out<=109;
				end
				if(in == 3) begin
					state<=6783;
					out<=110;
				end
				if(in == 4) begin
					state<=2894;
					out<=111;
				end
			end
			4784: begin
				if(in == 0) begin
					state<=4795;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=897;
					out<=114;
				end
				if(in == 3) begin
					state<=6784;
					out<=115;
				end
				if(in == 4) begin
					state<=2895;
					out<=116;
				end
			end
			4785: begin
				if(in == 0) begin
					state<=4796;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=898;
					out<=119;
				end
				if(in == 3) begin
					state<=6785;
					out<=120;
				end
				if(in == 4) begin
					state<=2896;
					out<=121;
				end
			end
			4786: begin
				if(in == 0) begin
					state<=4797;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=899;
					out<=124;
				end
				if(in == 3) begin
					state<=6786;
					out<=125;
				end
				if(in == 4) begin
					state<=2897;
					out<=126;
				end
			end
			4787: begin
				if(in == 0) begin
					state<=4788;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=890;
					out<=129;
				end
				if(in == 3) begin
					state<=6777;
					out<=130;
				end
				if(in == 4) begin
					state<=2888;
					out<=131;
				end
			end
			4788: begin
				if(in == 0) begin
					state<=4699;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=801;
					out<=134;
				end
				if(in == 3) begin
					state<=6688;
					out<=135;
				end
				if(in == 4) begin
					state<=2799;
					out<=136;
				end
			end
			4789: begin
				if(in == 0) begin
					state<=4700;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=802;
					out<=139;
				end
				if(in == 3) begin
					state<=6689;
					out<=140;
				end
				if(in == 4) begin
					state<=2800;
					out<=141;
				end
			end
			4790: begin
				if(in == 0) begin
					state<=4701;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=803;
					out<=144;
				end
				if(in == 3) begin
					state<=6690;
					out<=145;
				end
				if(in == 4) begin
					state<=2801;
					out<=146;
				end
			end
			4791: begin
				if(in == 0) begin
					state<=4702;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=804;
					out<=149;
				end
				if(in == 3) begin
					state<=6691;
					out<=150;
				end
				if(in == 4) begin
					state<=2802;
					out<=151;
				end
			end
			4792: begin
				if(in == 0) begin
					state<=4703;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=805;
					out<=154;
				end
				if(in == 3) begin
					state<=6692;
					out<=155;
				end
				if(in == 4) begin
					state<=2803;
					out<=156;
				end
			end
			4793: begin
				if(in == 0) begin
					state<=4704;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=806;
					out<=159;
				end
				if(in == 3) begin
					state<=6693;
					out<=160;
				end
				if(in == 4) begin
					state<=2804;
					out<=161;
				end
			end
			4794: begin
				if(in == 0) begin
					state<=4705;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=807;
					out<=164;
				end
				if(in == 3) begin
					state<=6694;
					out<=165;
				end
				if(in == 4) begin
					state<=2805;
					out<=166;
				end
			end
			4795: begin
				if(in == 0) begin
					state<=4706;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=808;
					out<=169;
				end
				if(in == 3) begin
					state<=6695;
					out<=170;
				end
				if(in == 4) begin
					state<=2806;
					out<=171;
				end
			end
			4796: begin
				if(in == 0) begin
					state<=4707;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=809;
					out<=174;
				end
				if(in == 3) begin
					state<=6696;
					out<=175;
				end
				if(in == 4) begin
					state<=2807;
					out<=176;
				end
			end
			4797: begin
				if(in == 0) begin
					state<=4698;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=800;
					out<=179;
				end
				if(in == 3) begin
					state<=6687;
					out<=180;
				end
				if(in == 4) begin
					state<=2798;
					out<=181;
				end
			end
			4798: begin
				if(in == 0) begin
					state<=4809;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=911;
					out<=184;
				end
				if(in == 3) begin
					state<=6176;
					out<=185;
				end
				if(in == 4) begin
					state<=2287;
					out<=186;
				end
			end
			4799: begin
				if(in == 0) begin
					state<=4810;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=912;
					out<=189;
				end
				if(in == 3) begin
					state<=6177;
					out<=190;
				end
				if(in == 4) begin
					state<=2288;
					out<=191;
				end
			end
			4800: begin
				if(in == 0) begin
					state<=4811;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=913;
					out<=194;
				end
				if(in == 3) begin
					state<=6178;
					out<=195;
				end
				if(in == 4) begin
					state<=2289;
					out<=196;
				end
			end
			4801: begin
				if(in == 0) begin
					state<=4812;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=914;
					out<=199;
				end
				if(in == 3) begin
					state<=6179;
					out<=200;
				end
				if(in == 4) begin
					state<=2290;
					out<=201;
				end
			end
			4802: begin
				if(in == 0) begin
					state<=4813;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=915;
					out<=204;
				end
				if(in == 3) begin
					state<=6180;
					out<=205;
				end
				if(in == 4) begin
					state<=2291;
					out<=206;
				end
			end
			4803: begin
				if(in == 0) begin
					state<=4814;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=916;
					out<=209;
				end
				if(in == 3) begin
					state<=6181;
					out<=210;
				end
				if(in == 4) begin
					state<=2292;
					out<=211;
				end
			end
			4804: begin
				if(in == 0) begin
					state<=4815;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=917;
					out<=214;
				end
				if(in == 3) begin
					state<=6182;
					out<=215;
				end
				if(in == 4) begin
					state<=2293;
					out<=216;
				end
			end
			4805: begin
				if(in == 0) begin
					state<=4816;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=918;
					out<=219;
				end
				if(in == 3) begin
					state<=6183;
					out<=220;
				end
				if(in == 4) begin
					state<=2294;
					out<=221;
				end
			end
			4806: begin
				if(in == 0) begin
					state<=4807;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=909;
					out<=224;
				end
				if(in == 3) begin
					state<=6174;
					out<=225;
				end
				if(in == 4) begin
					state<=2285;
					out<=226;
				end
			end
			4807: begin
				if(in == 0) begin
					state<=4818;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=920;
					out<=229;
				end
				if(in == 3) begin
					state<=6185;
					out<=230;
				end
				if(in == 4) begin
					state<=2296;
					out<=231;
				end
			end
			4808: begin
				if(in == 0) begin
					state<=4819;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=921;
					out<=234;
				end
				if(in == 3) begin
					state<=6186;
					out<=235;
				end
				if(in == 4) begin
					state<=2297;
					out<=236;
				end
			end
			4809: begin
				if(in == 0) begin
					state<=4820;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=922;
					out<=239;
				end
				if(in == 3) begin
					state<=6187;
					out<=240;
				end
				if(in == 4) begin
					state<=2298;
					out<=241;
				end
			end
			4810: begin
				if(in == 0) begin
					state<=4821;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=923;
					out<=244;
				end
				if(in == 3) begin
					state<=6188;
					out<=245;
				end
				if(in == 4) begin
					state<=2299;
					out<=246;
				end
			end
			4811: begin
				if(in == 0) begin
					state<=4822;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=924;
					out<=249;
				end
				if(in == 3) begin
					state<=6189;
					out<=250;
				end
				if(in == 4) begin
					state<=2300;
					out<=251;
				end
			end
			4812: begin
				if(in == 0) begin
					state<=4823;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=925;
					out<=254;
				end
				if(in == 3) begin
					state<=6190;
					out<=255;
				end
				if(in == 4) begin
					state<=2301;
					out<=0;
				end
			end
			4813: begin
				if(in == 0) begin
					state<=4824;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=926;
					out<=3;
				end
				if(in == 3) begin
					state<=6191;
					out<=4;
				end
				if(in == 4) begin
					state<=2302;
					out<=5;
				end
			end
			4814: begin
				if(in == 0) begin
					state<=4825;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=927;
					out<=8;
				end
				if(in == 3) begin
					state<=6192;
					out<=9;
				end
				if(in == 4) begin
					state<=2303;
					out<=10;
				end
			end
			4815: begin
				if(in == 0) begin
					state<=4826;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=928;
					out<=13;
				end
				if(in == 3) begin
					state<=6193;
					out<=14;
				end
				if(in == 4) begin
					state<=2304;
					out<=15;
				end
			end
			4816: begin
				if(in == 0) begin
					state<=4817;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=919;
					out<=18;
				end
				if(in == 3) begin
					state<=6184;
					out<=19;
				end
				if(in == 4) begin
					state<=2295;
					out<=20;
				end
			end
			4817: begin
				if(in == 0) begin
					state<=4828;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=930;
					out<=23;
				end
				if(in == 3) begin
					state<=6195;
					out<=24;
				end
				if(in == 4) begin
					state<=2306;
					out<=25;
				end
			end
			4818: begin
				if(in == 0) begin
					state<=4829;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=931;
					out<=28;
				end
				if(in == 3) begin
					state<=6196;
					out<=29;
				end
				if(in == 4) begin
					state<=2307;
					out<=30;
				end
			end
			4819: begin
				if(in == 0) begin
					state<=4830;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=932;
					out<=33;
				end
				if(in == 3) begin
					state<=6197;
					out<=34;
				end
				if(in == 4) begin
					state<=2308;
					out<=35;
				end
			end
			4820: begin
				if(in == 0) begin
					state<=4831;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=933;
					out<=38;
				end
				if(in == 3) begin
					state<=6198;
					out<=39;
				end
				if(in == 4) begin
					state<=2309;
					out<=40;
				end
			end
			4821: begin
				if(in == 0) begin
					state<=4832;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=934;
					out<=43;
				end
				if(in == 3) begin
					state<=6199;
					out<=44;
				end
				if(in == 4) begin
					state<=2310;
					out<=45;
				end
			end
			4822: begin
				if(in == 0) begin
					state<=4833;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=935;
					out<=48;
				end
				if(in == 3) begin
					state<=6200;
					out<=49;
				end
				if(in == 4) begin
					state<=2311;
					out<=50;
				end
			end
			4823: begin
				if(in == 0) begin
					state<=4834;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=936;
					out<=53;
				end
				if(in == 3) begin
					state<=6201;
					out<=54;
				end
				if(in == 4) begin
					state<=2312;
					out<=55;
				end
			end
			4824: begin
				if(in == 0) begin
					state<=4835;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=937;
					out<=58;
				end
				if(in == 3) begin
					state<=6202;
					out<=59;
				end
				if(in == 4) begin
					state<=2313;
					out<=60;
				end
			end
			4825: begin
				if(in == 0) begin
					state<=4836;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=938;
					out<=63;
				end
				if(in == 3) begin
					state<=6203;
					out<=64;
				end
				if(in == 4) begin
					state<=2314;
					out<=65;
				end
			end
			4826: begin
				if(in == 0) begin
					state<=4827;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=929;
					out<=68;
				end
				if(in == 3) begin
					state<=6194;
					out<=69;
				end
				if(in == 4) begin
					state<=2305;
					out<=70;
				end
			end
			4827: begin
				if(in == 0) begin
					state<=4838;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=940;
					out<=73;
				end
				if(in == 3) begin
					state<=6205;
					out<=74;
				end
				if(in == 4) begin
					state<=2316;
					out<=75;
				end
			end
			4828: begin
				if(in == 0) begin
					state<=4839;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=941;
					out<=78;
				end
				if(in == 3) begin
					state<=6206;
					out<=79;
				end
				if(in == 4) begin
					state<=2317;
					out<=80;
				end
			end
			4829: begin
				if(in == 0) begin
					state<=4840;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=942;
					out<=83;
				end
				if(in == 3) begin
					state<=6207;
					out<=84;
				end
				if(in == 4) begin
					state<=2318;
					out<=85;
				end
			end
			4830: begin
				if(in == 0) begin
					state<=4841;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=943;
					out<=88;
				end
				if(in == 3) begin
					state<=6208;
					out<=89;
				end
				if(in == 4) begin
					state<=2319;
					out<=90;
				end
			end
			4831: begin
				if(in == 0) begin
					state<=4842;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=944;
					out<=93;
				end
				if(in == 3) begin
					state<=6209;
					out<=94;
				end
				if(in == 4) begin
					state<=2320;
					out<=95;
				end
			end
			4832: begin
				if(in == 0) begin
					state<=4843;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=945;
					out<=98;
				end
				if(in == 3) begin
					state<=6210;
					out<=99;
				end
				if(in == 4) begin
					state<=2321;
					out<=100;
				end
			end
			4833: begin
				if(in == 0) begin
					state<=4844;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=946;
					out<=103;
				end
				if(in == 3) begin
					state<=6211;
					out<=104;
				end
				if(in == 4) begin
					state<=2322;
					out<=105;
				end
			end
			4834: begin
				if(in == 0) begin
					state<=4845;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=947;
					out<=108;
				end
				if(in == 3) begin
					state<=6212;
					out<=109;
				end
				if(in == 4) begin
					state<=2323;
					out<=110;
				end
			end
			4835: begin
				if(in == 0) begin
					state<=4846;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=948;
					out<=113;
				end
				if(in == 3) begin
					state<=6213;
					out<=114;
				end
				if(in == 4) begin
					state<=2324;
					out<=115;
				end
			end
			4836: begin
				if(in == 0) begin
					state<=4837;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=939;
					out<=118;
				end
				if(in == 3) begin
					state<=6204;
					out<=119;
				end
				if(in == 4) begin
					state<=2315;
					out<=120;
				end
			end
			4837: begin
				if(in == 0) begin
					state<=4848;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=950;
					out<=123;
				end
				if(in == 3) begin
					state<=6788;
					out<=124;
				end
				if(in == 4) begin
					state<=2899;
					out<=125;
				end
			end
			4838: begin
				if(in == 0) begin
					state<=4849;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=951;
					out<=128;
				end
				if(in == 3) begin
					state<=6789;
					out<=129;
				end
				if(in == 4) begin
					state<=2900;
					out<=130;
				end
			end
			4839: begin
				if(in == 0) begin
					state<=4850;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=952;
					out<=133;
				end
				if(in == 3) begin
					state<=6790;
					out<=134;
				end
				if(in == 4) begin
					state<=2901;
					out<=135;
				end
			end
			4840: begin
				if(in == 0) begin
					state<=4851;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=953;
					out<=138;
				end
				if(in == 3) begin
					state<=6791;
					out<=139;
				end
				if(in == 4) begin
					state<=2902;
					out<=140;
				end
			end
			4841: begin
				if(in == 0) begin
					state<=4852;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=954;
					out<=143;
				end
				if(in == 3) begin
					state<=6792;
					out<=144;
				end
				if(in == 4) begin
					state<=2903;
					out<=145;
				end
			end
			4842: begin
				if(in == 0) begin
					state<=4853;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=955;
					out<=148;
				end
				if(in == 3) begin
					state<=6793;
					out<=149;
				end
				if(in == 4) begin
					state<=2904;
					out<=150;
				end
			end
			4843: begin
				if(in == 0) begin
					state<=4854;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=956;
					out<=153;
				end
				if(in == 3) begin
					state<=6794;
					out<=154;
				end
				if(in == 4) begin
					state<=2905;
					out<=155;
				end
			end
			4844: begin
				if(in == 0) begin
					state<=4855;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=957;
					out<=158;
				end
				if(in == 3) begin
					state<=6795;
					out<=159;
				end
				if(in == 4) begin
					state<=2906;
					out<=160;
				end
			end
			4845: begin
				if(in == 0) begin
					state<=4856;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=958;
					out<=163;
				end
				if(in == 3) begin
					state<=6796;
					out<=164;
				end
				if(in == 4) begin
					state<=2907;
					out<=165;
				end
			end
			4846: begin
				if(in == 0) begin
					state<=4847;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=949;
					out<=168;
				end
				if(in == 3) begin
					state<=6787;
					out<=169;
				end
				if(in == 4) begin
					state<=2898;
					out<=170;
				end
			end
			4847: begin
				if(in == 0) begin
					state<=4858;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=960;
					out<=173;
				end
				if(in == 3) begin
					state<=6798;
					out<=174;
				end
				if(in == 4) begin
					state<=2909;
					out<=175;
				end
			end
			4848: begin
				if(in == 0) begin
					state<=4859;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=961;
					out<=178;
				end
				if(in == 3) begin
					state<=6799;
					out<=179;
				end
				if(in == 4) begin
					state<=2910;
					out<=180;
				end
			end
			4849: begin
				if(in == 0) begin
					state<=4860;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=962;
					out<=183;
				end
				if(in == 3) begin
					state<=6800;
					out<=184;
				end
				if(in == 4) begin
					state<=2911;
					out<=185;
				end
			end
			4850: begin
				if(in == 0) begin
					state<=4861;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=963;
					out<=188;
				end
				if(in == 3) begin
					state<=6801;
					out<=189;
				end
				if(in == 4) begin
					state<=2912;
					out<=190;
				end
			end
			4851: begin
				if(in == 0) begin
					state<=4862;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=964;
					out<=193;
				end
				if(in == 3) begin
					state<=6802;
					out<=194;
				end
				if(in == 4) begin
					state<=2913;
					out<=195;
				end
			end
			4852: begin
				if(in == 0) begin
					state<=4863;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=965;
					out<=198;
				end
				if(in == 3) begin
					state<=6803;
					out<=199;
				end
				if(in == 4) begin
					state<=2914;
					out<=200;
				end
			end
			4853: begin
				if(in == 0) begin
					state<=4864;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=966;
					out<=203;
				end
				if(in == 3) begin
					state<=6804;
					out<=204;
				end
				if(in == 4) begin
					state<=2915;
					out<=205;
				end
			end
			4854: begin
				if(in == 0) begin
					state<=4865;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=967;
					out<=208;
				end
				if(in == 3) begin
					state<=6805;
					out<=209;
				end
				if(in == 4) begin
					state<=2916;
					out<=210;
				end
			end
			4855: begin
				if(in == 0) begin
					state<=4866;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=968;
					out<=213;
				end
				if(in == 3) begin
					state<=6806;
					out<=214;
				end
				if(in == 4) begin
					state<=2917;
					out<=215;
				end
			end
			4856: begin
				if(in == 0) begin
					state<=4857;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=959;
					out<=218;
				end
				if(in == 3) begin
					state<=6797;
					out<=219;
				end
				if(in == 4) begin
					state<=2908;
					out<=220;
				end
			end
			4857: begin
				if(in == 0) begin
					state<=4868;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=970;
					out<=223;
				end
				if(in == 3) begin
					state<=6808;
					out<=224;
				end
				if(in == 4) begin
					state<=2919;
					out<=225;
				end
			end
			4858: begin
				if(in == 0) begin
					state<=4869;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=971;
					out<=228;
				end
				if(in == 3) begin
					state<=6809;
					out<=229;
				end
				if(in == 4) begin
					state<=2920;
					out<=230;
				end
			end
			4859: begin
				if(in == 0) begin
					state<=4870;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=972;
					out<=233;
				end
				if(in == 3) begin
					state<=6810;
					out<=234;
				end
				if(in == 4) begin
					state<=2921;
					out<=235;
				end
			end
			4860: begin
				if(in == 0) begin
					state<=4871;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=973;
					out<=238;
				end
				if(in == 3) begin
					state<=6811;
					out<=239;
				end
				if(in == 4) begin
					state<=2922;
					out<=240;
				end
			end
			4861: begin
				if(in == 0) begin
					state<=4872;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=974;
					out<=243;
				end
				if(in == 3) begin
					state<=6812;
					out<=244;
				end
				if(in == 4) begin
					state<=2923;
					out<=245;
				end
			end
			4862: begin
				if(in == 0) begin
					state<=4873;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=975;
					out<=248;
				end
				if(in == 3) begin
					state<=6813;
					out<=249;
				end
				if(in == 4) begin
					state<=2924;
					out<=250;
				end
			end
			4863: begin
				if(in == 0) begin
					state<=4874;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=976;
					out<=253;
				end
				if(in == 3) begin
					state<=6814;
					out<=254;
				end
				if(in == 4) begin
					state<=2925;
					out<=255;
				end
			end
			4864: begin
				if(in == 0) begin
					state<=4875;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=977;
					out<=2;
				end
				if(in == 3) begin
					state<=6815;
					out<=3;
				end
				if(in == 4) begin
					state<=2926;
					out<=4;
				end
			end
			4865: begin
				if(in == 0) begin
					state<=4876;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=978;
					out<=7;
				end
				if(in == 3) begin
					state<=6816;
					out<=8;
				end
				if(in == 4) begin
					state<=2927;
					out<=9;
				end
			end
			4866: begin
				if(in == 0) begin
					state<=4867;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=969;
					out<=12;
				end
				if(in == 3) begin
					state<=6807;
					out<=13;
				end
				if(in == 4) begin
					state<=2918;
					out<=14;
				end
			end
			4867: begin
				if(in == 0) begin
					state<=4878;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=980;
					out<=17;
				end
				if(in == 3) begin
					state<=6214;
					out<=18;
				end
				if(in == 4) begin
					state<=2325;
					out<=19;
				end
			end
			4868: begin
				if(in == 0) begin
					state<=4879;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=981;
					out<=22;
				end
				if(in == 3) begin
					state<=6215;
					out<=23;
				end
				if(in == 4) begin
					state<=2326;
					out<=24;
				end
			end
			4869: begin
				if(in == 0) begin
					state<=4880;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=982;
					out<=27;
				end
				if(in == 3) begin
					state<=6216;
					out<=28;
				end
				if(in == 4) begin
					state<=2327;
					out<=29;
				end
			end
			4870: begin
				if(in == 0) begin
					state<=4881;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=983;
					out<=32;
				end
				if(in == 3) begin
					state<=6217;
					out<=33;
				end
				if(in == 4) begin
					state<=2328;
					out<=34;
				end
			end
			4871: begin
				if(in == 0) begin
					state<=4882;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=984;
					out<=37;
				end
				if(in == 3) begin
					state<=6218;
					out<=38;
				end
				if(in == 4) begin
					state<=2329;
					out<=39;
				end
			end
			4872: begin
				if(in == 0) begin
					state<=4883;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=985;
					out<=42;
				end
				if(in == 3) begin
					state<=6219;
					out<=43;
				end
				if(in == 4) begin
					state<=2330;
					out<=44;
				end
			end
			4873: begin
				if(in == 0) begin
					state<=4884;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=986;
					out<=47;
				end
				if(in == 3) begin
					state<=6220;
					out<=48;
				end
				if(in == 4) begin
					state<=2331;
					out<=49;
				end
			end
			4874: begin
				if(in == 0) begin
					state<=4885;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=987;
					out<=52;
				end
				if(in == 3) begin
					state<=6221;
					out<=53;
				end
				if(in == 4) begin
					state<=2332;
					out<=54;
				end
			end
			4875: begin
				if(in == 0) begin
					state<=4886;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=988;
					out<=57;
				end
				if(in == 3) begin
					state<=6222;
					out<=58;
				end
				if(in == 4) begin
					state<=2333;
					out<=59;
				end
			end
			4876: begin
				if(in == 0) begin
					state<=4877;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=979;
					out<=62;
				end
				if(in == 3) begin
					state<=6817;
					out<=63;
				end
				if(in == 4) begin
					state<=2928;
					out<=64;
				end
			end
			4877: begin
				if(in == 0) begin
					state<=4888;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=990;
					out<=67;
				end
				if(in == 3) begin
					state<=6224;
					out<=68;
				end
				if(in == 4) begin
					state<=2335;
					out<=69;
				end
			end
			4878: begin
				if(in == 0) begin
					state<=4889;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=991;
					out<=72;
				end
				if(in == 3) begin
					state<=6225;
					out<=73;
				end
				if(in == 4) begin
					state<=2336;
					out<=74;
				end
			end
			4879: begin
				if(in == 0) begin
					state<=4890;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=992;
					out<=77;
				end
				if(in == 3) begin
					state<=6226;
					out<=78;
				end
				if(in == 4) begin
					state<=2337;
					out<=79;
				end
			end
			4880: begin
				if(in == 0) begin
					state<=4891;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=993;
					out<=82;
				end
				if(in == 3) begin
					state<=6227;
					out<=83;
				end
				if(in == 4) begin
					state<=2338;
					out<=84;
				end
			end
			4881: begin
				if(in == 0) begin
					state<=4892;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=994;
					out<=87;
				end
				if(in == 3) begin
					state<=6228;
					out<=88;
				end
				if(in == 4) begin
					state<=2339;
					out<=89;
				end
			end
			4882: begin
				if(in == 0) begin
					state<=4893;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=995;
					out<=92;
				end
				if(in == 3) begin
					state<=6229;
					out<=93;
				end
				if(in == 4) begin
					state<=2340;
					out<=94;
				end
			end
			4883: begin
				if(in == 0) begin
					state<=4894;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=996;
					out<=97;
				end
				if(in == 3) begin
					state<=6230;
					out<=98;
				end
				if(in == 4) begin
					state<=2341;
					out<=99;
				end
			end
			4884: begin
				if(in == 0) begin
					state<=4895;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=997;
					out<=102;
				end
				if(in == 3) begin
					state<=6231;
					out<=103;
				end
				if(in == 4) begin
					state<=2342;
					out<=104;
				end
			end
			4885: begin
				if(in == 0) begin
					state<=4896;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=998;
					out<=107;
				end
				if(in == 3) begin
					state<=6232;
					out<=108;
				end
				if(in == 4) begin
					state<=2343;
					out<=109;
				end
			end
			4886: begin
				if(in == 0) begin
					state<=4887;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=989;
					out<=112;
				end
				if(in == 3) begin
					state<=6223;
					out<=113;
				end
				if(in == 4) begin
					state<=2334;
					out<=114;
				end
			end
			4887: begin
				if(in == 0) begin
					state<=4245;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=347;
					out<=117;
				end
				if(in == 3) begin
					state<=6819;
					out<=118;
				end
				if(in == 4) begin
					state<=2930;
					out<=119;
				end
			end
			4888: begin
				if(in == 0) begin
					state<=4246;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=348;
					out<=122;
				end
				if(in == 3) begin
					state<=6820;
					out<=123;
				end
				if(in == 4) begin
					state<=2931;
					out<=124;
				end
			end
			4889: begin
				if(in == 0) begin
					state<=4247;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=349;
					out<=127;
				end
				if(in == 3) begin
					state<=6821;
					out<=128;
				end
				if(in == 4) begin
					state<=2932;
					out<=129;
				end
			end
			4890: begin
				if(in == 0) begin
					state<=4248;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=350;
					out<=132;
				end
				if(in == 3) begin
					state<=6822;
					out<=133;
				end
				if(in == 4) begin
					state<=2933;
					out<=134;
				end
			end
			4891: begin
				if(in == 0) begin
					state<=4249;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=351;
					out<=137;
				end
				if(in == 3) begin
					state<=6823;
					out<=138;
				end
				if(in == 4) begin
					state<=2934;
					out<=139;
				end
			end
			4892: begin
				if(in == 0) begin
					state<=4250;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=352;
					out<=142;
				end
				if(in == 3) begin
					state<=6824;
					out<=143;
				end
				if(in == 4) begin
					state<=2935;
					out<=144;
				end
			end
			4893: begin
				if(in == 0) begin
					state<=4251;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=353;
					out<=147;
				end
				if(in == 3) begin
					state<=6825;
					out<=148;
				end
				if(in == 4) begin
					state<=2936;
					out<=149;
				end
			end
			4894: begin
				if(in == 0) begin
					state<=4252;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=354;
					out<=152;
				end
				if(in == 3) begin
					state<=6826;
					out<=153;
				end
				if(in == 4) begin
					state<=2937;
					out<=154;
				end
			end
			4895: begin
				if(in == 0) begin
					state<=4253;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=355;
					out<=157;
				end
				if(in == 3) begin
					state<=6827;
					out<=158;
				end
				if(in == 4) begin
					state<=2938;
					out<=159;
				end
			end
			4896: begin
				if(in == 0) begin
					state<=4244;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=346;
					out<=162;
				end
				if(in == 3) begin
					state<=6818;
					out<=163;
				end
				if(in == 4) begin
					state<=2929;
					out<=164;
				end
			end
			4897: begin
				if(in == 0) begin
					state<=4908;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=1010;
					out<=167;
				end
				if(in == 3) begin
					state<=6879;
					out<=168;
				end
				if(in == 4) begin
					state<=2990;
					out<=169;
				end
			end
			4898: begin
				if(in == 0) begin
					state<=4909;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=1011;
					out<=172;
				end
				if(in == 3) begin
					state<=6880;
					out<=173;
				end
				if(in == 4) begin
					state<=2991;
					out<=174;
				end
			end
			4899: begin
				if(in == 0) begin
					state<=4910;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=1012;
					out<=177;
				end
				if(in == 3) begin
					state<=6881;
					out<=178;
				end
				if(in == 4) begin
					state<=2992;
					out<=179;
				end
			end
			4900: begin
				if(in == 0) begin
					state<=4911;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=1013;
					out<=182;
				end
				if(in == 3) begin
					state<=6882;
					out<=183;
				end
				if(in == 4) begin
					state<=2993;
					out<=184;
				end
			end
			4901: begin
				if(in == 0) begin
					state<=4912;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=1014;
					out<=187;
				end
				if(in == 3) begin
					state<=6883;
					out<=188;
				end
				if(in == 4) begin
					state<=2994;
					out<=189;
				end
			end
			4902: begin
				if(in == 0) begin
					state<=4913;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=1015;
					out<=192;
				end
				if(in == 3) begin
					state<=6884;
					out<=193;
				end
				if(in == 4) begin
					state<=2995;
					out<=194;
				end
			end
			4903: begin
				if(in == 0) begin
					state<=4914;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=1016;
					out<=197;
				end
				if(in == 3) begin
					state<=6885;
					out<=198;
				end
				if(in == 4) begin
					state<=2996;
					out<=199;
				end
			end
			4904: begin
				if(in == 0) begin
					state<=4915;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=1017;
					out<=202;
				end
				if(in == 3) begin
					state<=6886;
					out<=203;
				end
				if(in == 4) begin
					state<=2997;
					out<=204;
				end
			end
			4905: begin
				if(in == 0) begin
					state<=4916;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=1018;
					out<=207;
				end
				if(in == 3) begin
					state<=6887;
					out<=208;
				end
				if(in == 4) begin
					state<=2998;
					out<=209;
				end
			end
			4906: begin
				if(in == 0) begin
					state<=4907;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=1009;
					out<=212;
				end
				if(in == 3) begin
					state<=6878;
					out<=213;
				end
				if(in == 4) begin
					state<=2989;
					out<=214;
				end
			end
			4907: begin
				if(in == 0) begin
					state<=4918;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=1020;
					out<=217;
				end
				if(in == 3) begin
					state<=6889;
					out<=218;
				end
				if(in == 4) begin
					state<=3000;
					out<=219;
				end
			end
			4908: begin
				if(in == 0) begin
					state<=4919;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=1021;
					out<=222;
				end
				if(in == 3) begin
					state<=6890;
					out<=223;
				end
				if(in == 4) begin
					state<=3001;
					out<=224;
				end
			end
			4909: begin
				if(in == 0) begin
					state<=4920;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=1022;
					out<=227;
				end
				if(in == 3) begin
					state<=6891;
					out<=228;
				end
				if(in == 4) begin
					state<=3002;
					out<=229;
				end
			end
			4910: begin
				if(in == 0) begin
					state<=4921;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=1023;
					out<=232;
				end
				if(in == 3) begin
					state<=6892;
					out<=233;
				end
				if(in == 4) begin
					state<=3003;
					out<=234;
				end
			end
			4911: begin
				if(in == 0) begin
					state<=4922;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=1024;
					out<=237;
				end
				if(in == 3) begin
					state<=6893;
					out<=238;
				end
				if(in == 4) begin
					state<=3004;
					out<=239;
				end
			end
			4912: begin
				if(in == 0) begin
					state<=4923;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=1025;
					out<=242;
				end
				if(in == 3) begin
					state<=6894;
					out<=243;
				end
				if(in == 4) begin
					state<=3005;
					out<=244;
				end
			end
			4913: begin
				if(in == 0) begin
					state<=4924;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=1026;
					out<=247;
				end
				if(in == 3) begin
					state<=6895;
					out<=248;
				end
				if(in == 4) begin
					state<=3006;
					out<=249;
				end
			end
			4914: begin
				if(in == 0) begin
					state<=4925;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=1027;
					out<=252;
				end
				if(in == 3) begin
					state<=6896;
					out<=253;
				end
				if(in == 4) begin
					state<=3007;
					out<=254;
				end
			end
			4915: begin
				if(in == 0) begin
					state<=4926;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=1028;
					out<=1;
				end
				if(in == 3) begin
					state<=6897;
					out<=2;
				end
				if(in == 4) begin
					state<=3008;
					out<=3;
				end
			end
			4916: begin
				if(in == 0) begin
					state<=4917;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=1019;
					out<=6;
				end
				if(in == 3) begin
					state<=6888;
					out<=7;
				end
				if(in == 4) begin
					state<=2999;
					out<=8;
				end
			end
			4917: begin
				if(in == 0) begin
					state<=4294;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=396;
					out<=11;
				end
				if(in == 3) begin
					state<=6899;
					out<=12;
				end
				if(in == 4) begin
					state<=3010;
					out<=13;
				end
			end
			4918: begin
				if(in == 0) begin
					state<=4295;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=397;
					out<=16;
				end
				if(in == 3) begin
					state<=6900;
					out<=17;
				end
				if(in == 4) begin
					state<=3011;
					out<=18;
				end
			end
			4919: begin
				if(in == 0) begin
					state<=4296;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=398;
					out<=21;
				end
				if(in == 3) begin
					state<=6901;
					out<=22;
				end
				if(in == 4) begin
					state<=3012;
					out<=23;
				end
			end
			4920: begin
				if(in == 0) begin
					state<=4297;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=399;
					out<=26;
				end
				if(in == 3) begin
					state<=6902;
					out<=27;
				end
				if(in == 4) begin
					state<=3013;
					out<=28;
				end
			end
			4921: begin
				if(in == 0) begin
					state<=4298;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=400;
					out<=31;
				end
				if(in == 3) begin
					state<=6903;
					out<=32;
				end
				if(in == 4) begin
					state<=3014;
					out<=33;
				end
			end
			4922: begin
				if(in == 0) begin
					state<=4299;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=401;
					out<=36;
				end
				if(in == 3) begin
					state<=6904;
					out<=37;
				end
				if(in == 4) begin
					state<=3015;
					out<=38;
				end
			end
			4923: begin
				if(in == 0) begin
					state<=4300;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=402;
					out<=41;
				end
				if(in == 3) begin
					state<=6905;
					out<=42;
				end
				if(in == 4) begin
					state<=3016;
					out<=43;
				end
			end
			4924: begin
				if(in == 0) begin
					state<=4301;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=403;
					out<=46;
				end
				if(in == 3) begin
					state<=6906;
					out<=47;
				end
				if(in == 4) begin
					state<=3017;
					out<=48;
				end
			end
			4925: begin
				if(in == 0) begin
					state<=4302;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=404;
					out<=51;
				end
				if(in == 3) begin
					state<=6907;
					out<=52;
				end
				if(in == 4) begin
					state<=3018;
					out<=53;
				end
			end
			4926: begin
				if(in == 0) begin
					state<=4927;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=1029;
					out<=56;
				end
				if(in == 3) begin
					state<=6898;
					out<=57;
				end
				if(in == 4) begin
					state<=3009;
					out<=58;
				end
			end
			4927: begin
				if(in == 0) begin
					state<=4304;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=406;
					out<=61;
				end
				if(in == 3) begin
					state<=6909;
					out<=62;
				end
				if(in == 4) begin
					state<=3020;
					out<=63;
				end
			end
			4928: begin
				if(in == 0) begin
					state<=4939;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=1041;
					out<=66;
				end
				if(in == 3) begin
					state<=6929;
					out<=67;
				end
				if(in == 4) begin
					state<=3040;
					out<=68;
				end
			end
			4929: begin
				if(in == 0) begin
					state<=4940;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=1042;
					out<=71;
				end
				if(in == 3) begin
					state<=6930;
					out<=72;
				end
				if(in == 4) begin
					state<=3041;
					out<=73;
				end
			end
			4930: begin
				if(in == 0) begin
					state<=4941;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=1043;
					out<=76;
				end
				if(in == 3) begin
					state<=6931;
					out<=77;
				end
				if(in == 4) begin
					state<=3042;
					out<=78;
				end
			end
			4931: begin
				if(in == 0) begin
					state<=4942;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=1044;
					out<=81;
				end
				if(in == 3) begin
					state<=6932;
					out<=82;
				end
				if(in == 4) begin
					state<=3043;
					out<=83;
				end
			end
			4932: begin
				if(in == 0) begin
					state<=4943;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=1045;
					out<=86;
				end
				if(in == 3) begin
					state<=6933;
					out<=87;
				end
				if(in == 4) begin
					state<=3044;
					out<=88;
				end
			end
			4933: begin
				if(in == 0) begin
					state<=4944;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=1046;
					out<=91;
				end
				if(in == 3) begin
					state<=6934;
					out<=92;
				end
				if(in == 4) begin
					state<=3045;
					out<=93;
				end
			end
			4934: begin
				if(in == 0) begin
					state<=4945;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=1047;
					out<=96;
				end
				if(in == 3) begin
					state<=6935;
					out<=97;
				end
				if(in == 4) begin
					state<=3046;
					out<=98;
				end
			end
			4935: begin
				if(in == 0) begin
					state<=4946;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=1048;
					out<=101;
				end
				if(in == 3) begin
					state<=6936;
					out<=102;
				end
				if(in == 4) begin
					state<=3047;
					out<=103;
				end
			end
			4936: begin
				if(in == 0) begin
					state<=4947;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=1049;
					out<=106;
				end
				if(in == 3) begin
					state<=6937;
					out<=107;
				end
				if(in == 4) begin
					state<=3048;
					out<=108;
				end
			end
			4937: begin
				if(in == 0) begin
					state<=4938;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=1040;
					out<=111;
				end
				if(in == 3) begin
					state<=6928;
					out<=112;
				end
				if(in == 4) begin
					state<=3039;
					out<=113;
				end
			end
			4938: begin
				if(in == 0) begin
					state<=4949;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=1051;
					out<=116;
				end
				if(in == 3) begin
					state<=6939;
					out<=117;
				end
				if(in == 4) begin
					state<=3050;
					out<=118;
				end
			end
			4939: begin
				if(in == 0) begin
					state<=4950;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=1052;
					out<=121;
				end
				if(in == 3) begin
					state<=6940;
					out<=122;
				end
				if(in == 4) begin
					state<=3051;
					out<=123;
				end
			end
			4940: begin
				if(in == 0) begin
					state<=4951;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=1053;
					out<=126;
				end
				if(in == 3) begin
					state<=6941;
					out<=127;
				end
				if(in == 4) begin
					state<=3052;
					out<=128;
				end
			end
			4941: begin
				if(in == 0) begin
					state<=4952;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=1054;
					out<=131;
				end
				if(in == 3) begin
					state<=6942;
					out<=132;
				end
				if(in == 4) begin
					state<=3053;
					out<=133;
				end
			end
			4942: begin
				if(in == 0) begin
					state<=4953;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=1055;
					out<=136;
				end
				if(in == 3) begin
					state<=6943;
					out<=137;
				end
				if(in == 4) begin
					state<=3054;
					out<=138;
				end
			end
			4943: begin
				if(in == 0) begin
					state<=4954;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=1056;
					out<=141;
				end
				if(in == 3) begin
					state<=6944;
					out<=142;
				end
				if(in == 4) begin
					state<=3055;
					out<=143;
				end
			end
			4944: begin
				if(in == 0) begin
					state<=4955;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=1057;
					out<=146;
				end
				if(in == 3) begin
					state<=6945;
					out<=147;
				end
				if(in == 4) begin
					state<=3056;
					out<=148;
				end
			end
			4945: begin
				if(in == 0) begin
					state<=4956;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=1058;
					out<=151;
				end
				if(in == 3) begin
					state<=6946;
					out<=152;
				end
				if(in == 4) begin
					state<=3057;
					out<=153;
				end
			end
			4946: begin
				if(in == 0) begin
					state<=4957;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=1059;
					out<=156;
				end
				if(in == 3) begin
					state<=6947;
					out<=157;
				end
				if(in == 4) begin
					state<=3058;
					out<=158;
				end
			end
			4947: begin
				if(in == 0) begin
					state<=4948;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=1050;
					out<=161;
				end
				if(in == 3) begin
					state<=6938;
					out<=162;
				end
				if(in == 4) begin
					state<=3049;
					out<=163;
				end
			end
			4948: begin
				if(in == 0) begin
					state<=4959;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=1061;
					out<=166;
				end
				if(in == 3) begin
					state<=6949;
					out<=167;
				end
				if(in == 4) begin
					state<=3060;
					out<=168;
				end
			end
			4949: begin
				if(in == 0) begin
					state<=4960;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=1062;
					out<=171;
				end
				if(in == 3) begin
					state<=6950;
					out<=172;
				end
				if(in == 4) begin
					state<=3061;
					out<=173;
				end
			end
			4950: begin
				if(in == 0) begin
					state<=4961;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=1063;
					out<=176;
				end
				if(in == 3) begin
					state<=6951;
					out<=177;
				end
				if(in == 4) begin
					state<=3062;
					out<=178;
				end
			end
			4951: begin
				if(in == 0) begin
					state<=4962;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=1064;
					out<=181;
				end
				if(in == 3) begin
					state<=6952;
					out<=182;
				end
				if(in == 4) begin
					state<=3063;
					out<=183;
				end
			end
			4952: begin
				if(in == 0) begin
					state<=4963;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=1065;
					out<=186;
				end
				if(in == 3) begin
					state<=6953;
					out<=187;
				end
				if(in == 4) begin
					state<=3064;
					out<=188;
				end
			end
			4953: begin
				if(in == 0) begin
					state<=4964;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=1066;
					out<=191;
				end
				if(in == 3) begin
					state<=6954;
					out<=192;
				end
				if(in == 4) begin
					state<=3065;
					out<=193;
				end
			end
			4954: begin
				if(in == 0) begin
					state<=4965;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=1067;
					out<=196;
				end
				if(in == 3) begin
					state<=6955;
					out<=197;
				end
				if(in == 4) begin
					state<=3066;
					out<=198;
				end
			end
			4955: begin
				if(in == 0) begin
					state<=4966;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=1068;
					out<=201;
				end
				if(in == 3) begin
					state<=6956;
					out<=202;
				end
				if(in == 4) begin
					state<=3067;
					out<=203;
				end
			end
			4956: begin
				if(in == 0) begin
					state<=4967;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=1069;
					out<=206;
				end
				if(in == 3) begin
					state<=6957;
					out<=207;
				end
				if(in == 4) begin
					state<=3068;
					out<=208;
				end
			end
			4957: begin
				if(in == 0) begin
					state<=4958;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=1060;
					out<=211;
				end
				if(in == 3) begin
					state<=6948;
					out<=212;
				end
				if(in == 4) begin
					state<=3059;
					out<=213;
				end
			end
			4958: begin
				if(in == 0) begin
					state<=4969;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=1071;
					out<=216;
				end
				if(in == 3) begin
					state<=6959;
					out<=217;
				end
				if(in == 4) begin
					state<=3070;
					out<=218;
				end
			end
			4959: begin
				if(in == 0) begin
					state<=4970;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=1072;
					out<=221;
				end
				if(in == 3) begin
					state<=6960;
					out<=222;
				end
				if(in == 4) begin
					state<=3071;
					out<=223;
				end
			end
			4960: begin
				if(in == 0) begin
					state<=4971;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=1073;
					out<=226;
				end
				if(in == 3) begin
					state<=6961;
					out<=227;
				end
				if(in == 4) begin
					state<=3072;
					out<=228;
				end
			end
			4961: begin
				if(in == 0) begin
					state<=4972;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=1074;
					out<=231;
				end
				if(in == 3) begin
					state<=6962;
					out<=232;
				end
				if(in == 4) begin
					state<=3073;
					out<=233;
				end
			end
			4962: begin
				if(in == 0) begin
					state<=4973;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=1075;
					out<=236;
				end
				if(in == 3) begin
					state<=6963;
					out<=237;
				end
				if(in == 4) begin
					state<=3074;
					out<=238;
				end
			end
			4963: begin
				if(in == 0) begin
					state<=4974;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=1076;
					out<=241;
				end
				if(in == 3) begin
					state<=6964;
					out<=242;
				end
				if(in == 4) begin
					state<=3075;
					out<=243;
				end
			end
			4964: begin
				if(in == 0) begin
					state<=4975;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=1077;
					out<=246;
				end
				if(in == 3) begin
					state<=6965;
					out<=247;
				end
				if(in == 4) begin
					state<=3076;
					out<=248;
				end
			end
			4965: begin
				if(in == 0) begin
					state<=4976;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=1078;
					out<=251;
				end
				if(in == 3) begin
					state<=6966;
					out<=252;
				end
				if(in == 4) begin
					state<=3077;
					out<=253;
				end
			end
			4966: begin
				if(in == 0) begin
					state<=4977;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=1079;
					out<=0;
				end
				if(in == 3) begin
					state<=6967;
					out<=1;
				end
				if(in == 4) begin
					state<=3078;
					out<=2;
				end
			end
			4967: begin
				if(in == 0) begin
					state<=4968;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=1070;
					out<=5;
				end
				if(in == 3) begin
					state<=6958;
					out<=6;
				end
				if(in == 4) begin
					state<=3069;
					out<=7;
				end
			end
			4968: begin
				if(in == 0) begin
					state<=4979;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=1081;
					out<=10;
				end
				if(in == 3) begin
					state<=6969;
					out<=11;
				end
				if(in == 4) begin
					state<=3080;
					out<=12;
				end
			end
			4969: begin
				if(in == 0) begin
					state<=4980;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=1082;
					out<=15;
				end
				if(in == 3) begin
					state<=6970;
					out<=16;
				end
				if(in == 4) begin
					state<=3081;
					out<=17;
				end
			end
			4970: begin
				if(in == 0) begin
					state<=4981;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=1083;
					out<=20;
				end
				if(in == 3) begin
					state<=6971;
					out<=21;
				end
				if(in == 4) begin
					state<=3082;
					out<=22;
				end
			end
			4971: begin
				if(in == 0) begin
					state<=4982;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=1084;
					out<=25;
				end
				if(in == 3) begin
					state<=6972;
					out<=26;
				end
				if(in == 4) begin
					state<=3083;
					out<=27;
				end
			end
			4972: begin
				if(in == 0) begin
					state<=4983;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=1085;
					out<=30;
				end
				if(in == 3) begin
					state<=6973;
					out<=31;
				end
				if(in == 4) begin
					state<=3084;
					out<=32;
				end
			end
			4973: begin
				if(in == 0) begin
					state<=4984;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=1086;
					out<=35;
				end
				if(in == 3) begin
					state<=6974;
					out<=36;
				end
				if(in == 4) begin
					state<=3085;
					out<=37;
				end
			end
			4974: begin
				if(in == 0) begin
					state<=4985;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=1087;
					out<=40;
				end
				if(in == 3) begin
					state<=6975;
					out<=41;
				end
				if(in == 4) begin
					state<=3086;
					out<=42;
				end
			end
			4975: begin
				if(in == 0) begin
					state<=4986;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=1088;
					out<=45;
				end
				if(in == 3) begin
					state<=6976;
					out<=46;
				end
				if(in == 4) begin
					state<=3087;
					out<=47;
				end
			end
			4976: begin
				if(in == 0) begin
					state<=4987;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=1089;
					out<=50;
				end
				if(in == 3) begin
					state<=6977;
					out<=51;
				end
				if(in == 4) begin
					state<=3088;
					out<=52;
				end
			end
			4977: begin
				if(in == 0) begin
					state<=4978;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=1080;
					out<=55;
				end
				if(in == 3) begin
					state<=6968;
					out<=56;
				end
				if(in == 4) begin
					state<=3079;
					out<=57;
				end
			end
			4978: begin
				if(in == 0) begin
					state<=4989;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=1091;
					out<=60;
				end
				if(in == 3) begin
					state<=6979;
					out<=61;
				end
				if(in == 4) begin
					state<=3090;
					out<=62;
				end
			end
			4979: begin
				if(in == 0) begin
					state<=4990;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=1092;
					out<=65;
				end
				if(in == 3) begin
					state<=6980;
					out<=66;
				end
				if(in == 4) begin
					state<=3091;
					out<=67;
				end
			end
			4980: begin
				if(in == 0) begin
					state<=4991;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=1093;
					out<=70;
				end
				if(in == 3) begin
					state<=6981;
					out<=71;
				end
				if(in == 4) begin
					state<=3092;
					out<=72;
				end
			end
			4981: begin
				if(in == 0) begin
					state<=4992;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=1094;
					out<=75;
				end
				if(in == 3) begin
					state<=6982;
					out<=76;
				end
				if(in == 4) begin
					state<=3093;
					out<=77;
				end
			end
			4982: begin
				if(in == 0) begin
					state<=4993;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=1095;
					out<=80;
				end
				if(in == 3) begin
					state<=6983;
					out<=81;
				end
				if(in == 4) begin
					state<=3094;
					out<=82;
				end
			end
			4983: begin
				if(in == 0) begin
					state<=4994;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=1096;
					out<=85;
				end
				if(in == 3) begin
					state<=6984;
					out<=86;
				end
				if(in == 4) begin
					state<=3095;
					out<=87;
				end
			end
			4984: begin
				if(in == 0) begin
					state<=4995;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=1097;
					out<=90;
				end
				if(in == 3) begin
					state<=6985;
					out<=91;
				end
				if(in == 4) begin
					state<=3096;
					out<=92;
				end
			end
			4985: begin
				if(in == 0) begin
					state<=4996;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=1098;
					out<=95;
				end
				if(in == 3) begin
					state<=6986;
					out<=96;
				end
				if(in == 4) begin
					state<=3097;
					out<=97;
				end
			end
			4986: begin
				if(in == 0) begin
					state<=4997;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=1099;
					out<=100;
				end
				if(in == 3) begin
					state<=6987;
					out<=101;
				end
				if(in == 4) begin
					state<=3098;
					out<=102;
				end
			end
			4987: begin
				if(in == 0) begin
					state<=4988;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=1090;
					out<=105;
				end
				if(in == 3) begin
					state<=6978;
					out<=106;
				end
				if(in == 4) begin
					state<=3089;
					out<=107;
				end
			end
			4988: begin
				if(in == 0) begin
					state<=4999;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=1101;
					out<=110;
				end
				if(in == 3) begin
					state<=6989;
					out<=111;
				end
				if(in == 4) begin
					state<=3100;
					out<=112;
				end
			end
			4989: begin
				if(in == 0) begin
					state<=5000;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=1102;
					out<=115;
				end
				if(in == 3) begin
					state<=6990;
					out<=116;
				end
				if(in == 4) begin
					state<=3101;
					out<=117;
				end
			end
			4990: begin
				if(in == 0) begin
					state<=5001;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=1103;
					out<=120;
				end
				if(in == 3) begin
					state<=6991;
					out<=121;
				end
				if(in == 4) begin
					state<=3102;
					out<=122;
				end
			end
			4991: begin
				if(in == 0) begin
					state<=5002;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=1104;
					out<=125;
				end
				if(in == 3) begin
					state<=6992;
					out<=126;
				end
				if(in == 4) begin
					state<=3103;
					out<=127;
				end
			end
			4992: begin
				if(in == 0) begin
					state<=5003;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=1105;
					out<=130;
				end
				if(in == 3) begin
					state<=6993;
					out<=131;
				end
				if(in == 4) begin
					state<=3104;
					out<=132;
				end
			end
			4993: begin
				if(in == 0) begin
					state<=5004;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=1106;
					out<=135;
				end
				if(in == 3) begin
					state<=6994;
					out<=136;
				end
				if(in == 4) begin
					state<=3105;
					out<=137;
				end
			end
			4994: begin
				if(in == 0) begin
					state<=5005;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=1107;
					out<=140;
				end
				if(in == 3) begin
					state<=6995;
					out<=141;
				end
				if(in == 4) begin
					state<=3106;
					out<=142;
				end
			end
			4995: begin
				if(in == 0) begin
					state<=5006;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=1108;
					out<=145;
				end
				if(in == 3) begin
					state<=6996;
					out<=146;
				end
				if(in == 4) begin
					state<=3107;
					out<=147;
				end
			end
			4996: begin
				if(in == 0) begin
					state<=5007;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=1109;
					out<=150;
				end
				if(in == 3) begin
					state<=6997;
					out<=151;
				end
				if(in == 4) begin
					state<=3108;
					out<=152;
				end
			end
			4997: begin
				if(in == 0) begin
					state<=4998;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=1100;
					out<=155;
				end
				if(in == 3) begin
					state<=6988;
					out<=156;
				end
				if(in == 4) begin
					state<=3099;
					out<=157;
				end
			end
			4998: begin
				if(in == 0) begin
					state<=5009;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=1111;
					out<=160;
				end
				if(in == 3) begin
					state<=6999;
					out<=161;
				end
				if(in == 4) begin
					state<=3110;
					out<=162;
				end
			end
			4999: begin
				if(in == 0) begin
					state<=5010;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=1112;
					out<=165;
				end
				if(in == 3) begin
					state<=7000;
					out<=166;
				end
				if(in == 4) begin
					state<=3111;
					out<=167;
				end
			end
			5000: begin
				if(in == 0) begin
					state<=5011;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=1113;
					out<=170;
				end
				if(in == 3) begin
					state<=7001;
					out<=171;
				end
				if(in == 4) begin
					state<=3112;
					out<=172;
				end
			end
			5001: begin
				if(in == 0) begin
					state<=5012;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=1114;
					out<=175;
				end
				if(in == 3) begin
					state<=7002;
					out<=176;
				end
				if(in == 4) begin
					state<=3113;
					out<=177;
				end
			end
			5002: begin
				if(in == 0) begin
					state<=5013;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=1115;
					out<=180;
				end
				if(in == 3) begin
					state<=7003;
					out<=181;
				end
				if(in == 4) begin
					state<=3114;
					out<=182;
				end
			end
			5003: begin
				if(in == 0) begin
					state<=5014;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=1116;
					out<=185;
				end
				if(in == 3) begin
					state<=7004;
					out<=186;
				end
				if(in == 4) begin
					state<=3115;
					out<=187;
				end
			end
			5004: begin
				if(in == 0) begin
					state<=5015;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=1117;
					out<=190;
				end
				if(in == 3) begin
					state<=7005;
					out<=191;
				end
				if(in == 4) begin
					state<=3116;
					out<=192;
				end
			end
			5005: begin
				if(in == 0) begin
					state<=5016;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=1118;
					out<=195;
				end
				if(in == 3) begin
					state<=7006;
					out<=196;
				end
				if(in == 4) begin
					state<=3117;
					out<=197;
				end
			end
			5006: begin
				if(in == 0) begin
					state<=5017;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=1119;
					out<=200;
				end
				if(in == 3) begin
					state<=7007;
					out<=201;
				end
				if(in == 4) begin
					state<=3118;
					out<=202;
				end
			end
			5007: begin
				if(in == 0) begin
					state<=5008;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=1110;
					out<=205;
				end
				if(in == 3) begin
					state<=6998;
					out<=206;
				end
				if(in == 4) begin
					state<=3109;
					out<=207;
				end
			end
			5008: begin
				if(in == 0) begin
					state<=5019;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=1121;
					out<=210;
				end
				if(in == 3) begin
					state<=7009;
					out<=211;
				end
				if(in == 4) begin
					state<=3120;
					out<=212;
				end
			end
			5009: begin
				if(in == 0) begin
					state<=5020;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=1122;
					out<=215;
				end
				if(in == 3) begin
					state<=7010;
					out<=216;
				end
				if(in == 4) begin
					state<=3121;
					out<=217;
				end
			end
			5010: begin
				if(in == 0) begin
					state<=5021;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=1123;
					out<=220;
				end
				if(in == 3) begin
					state<=7011;
					out<=221;
				end
				if(in == 4) begin
					state<=3122;
					out<=222;
				end
			end
			5011: begin
				if(in == 0) begin
					state<=5022;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=1124;
					out<=225;
				end
				if(in == 3) begin
					state<=7012;
					out<=226;
				end
				if(in == 4) begin
					state<=3123;
					out<=227;
				end
			end
			5012: begin
				if(in == 0) begin
					state<=5023;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=1125;
					out<=230;
				end
				if(in == 3) begin
					state<=7013;
					out<=231;
				end
				if(in == 4) begin
					state<=3124;
					out<=232;
				end
			end
			5013: begin
				if(in == 0) begin
					state<=5024;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=1126;
					out<=235;
				end
				if(in == 3) begin
					state<=7014;
					out<=236;
				end
				if(in == 4) begin
					state<=3125;
					out<=237;
				end
			end
			5014: begin
				if(in == 0) begin
					state<=5025;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=1127;
					out<=240;
				end
				if(in == 3) begin
					state<=7015;
					out<=241;
				end
				if(in == 4) begin
					state<=3126;
					out<=242;
				end
			end
			5015: begin
				if(in == 0) begin
					state<=5026;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=1128;
					out<=245;
				end
				if(in == 3) begin
					state<=7016;
					out<=246;
				end
				if(in == 4) begin
					state<=3127;
					out<=247;
				end
			end
			5016: begin
				if(in == 0) begin
					state<=5027;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=1129;
					out<=250;
				end
				if(in == 3) begin
					state<=7017;
					out<=251;
				end
				if(in == 4) begin
					state<=3128;
					out<=252;
				end
			end
			5017: begin
				if(in == 0) begin
					state<=5018;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=1120;
					out<=255;
				end
				if(in == 3) begin
					state<=7008;
					out<=0;
				end
				if(in == 4) begin
					state<=3119;
					out<=1;
				end
			end
			5018: begin
				if(in == 0) begin
					state<=5029;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=1131;
					out<=4;
				end
				if(in == 3) begin
					state<=7019;
					out<=5;
				end
				if(in == 4) begin
					state<=3130;
					out<=6;
				end
			end
			5019: begin
				if(in == 0) begin
					state<=5030;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=1132;
					out<=9;
				end
				if(in == 3) begin
					state<=7020;
					out<=10;
				end
				if(in == 4) begin
					state<=3131;
					out<=11;
				end
			end
			5020: begin
				if(in == 0) begin
					state<=5031;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=1133;
					out<=14;
				end
				if(in == 3) begin
					state<=7021;
					out<=15;
				end
				if(in == 4) begin
					state<=3132;
					out<=16;
				end
			end
			5021: begin
				if(in == 0) begin
					state<=5032;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=1134;
					out<=19;
				end
				if(in == 3) begin
					state<=7022;
					out<=20;
				end
				if(in == 4) begin
					state<=3133;
					out<=21;
				end
			end
			5022: begin
				if(in == 0) begin
					state<=5033;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=1135;
					out<=24;
				end
				if(in == 3) begin
					state<=7023;
					out<=25;
				end
				if(in == 4) begin
					state<=3134;
					out<=26;
				end
			end
			5023: begin
				if(in == 0) begin
					state<=5034;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=1136;
					out<=29;
				end
				if(in == 3) begin
					state<=7024;
					out<=30;
				end
				if(in == 4) begin
					state<=3135;
					out<=31;
				end
			end
			5024: begin
				if(in == 0) begin
					state<=5035;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=1137;
					out<=34;
				end
				if(in == 3) begin
					state<=7025;
					out<=35;
				end
				if(in == 4) begin
					state<=3136;
					out<=36;
				end
			end
			5025: begin
				if(in == 0) begin
					state<=5036;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=1138;
					out<=39;
				end
				if(in == 3) begin
					state<=7026;
					out<=40;
				end
				if(in == 4) begin
					state<=3137;
					out<=41;
				end
			end
			5026: begin
				if(in == 0) begin
					state<=5037;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=1139;
					out<=44;
				end
				if(in == 3) begin
					state<=7027;
					out<=45;
				end
				if(in == 4) begin
					state<=3138;
					out<=46;
				end
			end
			5027: begin
				if(in == 0) begin
					state<=5028;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=1130;
					out<=49;
				end
				if(in == 3) begin
					state<=7018;
					out<=50;
				end
				if(in == 4) begin
					state<=3129;
					out<=51;
				end
			end
			5028: begin
				if(in == 0) begin
					state<=5039;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=1141;
					out<=54;
				end
				if(in == 3) begin
					state<=7029;
					out<=55;
				end
				if(in == 4) begin
					state<=3140;
					out<=56;
				end
			end
			5029: begin
				if(in == 0) begin
					state<=5040;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=1142;
					out<=59;
				end
				if(in == 3) begin
					state<=7030;
					out<=60;
				end
				if(in == 4) begin
					state<=3141;
					out<=61;
				end
			end
			5030: begin
				if(in == 0) begin
					state<=5041;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=1143;
					out<=64;
				end
				if(in == 3) begin
					state<=7031;
					out<=65;
				end
				if(in == 4) begin
					state<=3142;
					out<=66;
				end
			end
			5031: begin
				if(in == 0) begin
					state<=5042;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=1144;
					out<=69;
				end
				if(in == 3) begin
					state<=7032;
					out<=70;
				end
				if(in == 4) begin
					state<=3143;
					out<=71;
				end
			end
			5032: begin
				if(in == 0) begin
					state<=5043;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=1145;
					out<=74;
				end
				if(in == 3) begin
					state<=7033;
					out<=75;
				end
				if(in == 4) begin
					state<=3144;
					out<=76;
				end
			end
			5033: begin
				if(in == 0) begin
					state<=5044;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=1146;
					out<=79;
				end
				if(in == 3) begin
					state<=7034;
					out<=80;
				end
				if(in == 4) begin
					state<=3145;
					out<=81;
				end
			end
			5034: begin
				if(in == 0) begin
					state<=5045;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=1147;
					out<=84;
				end
				if(in == 3) begin
					state<=7035;
					out<=85;
				end
				if(in == 4) begin
					state<=3146;
					out<=86;
				end
			end
			5035: begin
				if(in == 0) begin
					state<=5046;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=1148;
					out<=89;
				end
				if(in == 3) begin
					state<=7036;
					out<=90;
				end
				if(in == 4) begin
					state<=3147;
					out<=91;
				end
			end
			5036: begin
				if(in == 0) begin
					state<=5047;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=1149;
					out<=94;
				end
				if(in == 3) begin
					state<=7037;
					out<=95;
				end
				if(in == 4) begin
					state<=3148;
					out<=96;
				end
			end
			5037: begin
				if(in == 0) begin
					state<=5038;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=1140;
					out<=99;
				end
				if(in == 3) begin
					state<=7028;
					out<=100;
				end
				if(in == 4) begin
					state<=3139;
					out<=101;
				end
			end
			5038: begin
				if(in == 0) begin
					state<=5049;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=1151;
					out<=104;
				end
				if(in == 3) begin
					state<=7039;
					out<=105;
				end
				if(in == 4) begin
					state<=3150;
					out<=106;
				end
			end
			5039: begin
				if(in == 0) begin
					state<=5050;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=1152;
					out<=109;
				end
				if(in == 3) begin
					state<=7040;
					out<=110;
				end
				if(in == 4) begin
					state<=3151;
					out<=111;
				end
			end
			5040: begin
				if(in == 0) begin
					state<=5051;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=1153;
					out<=114;
				end
				if(in == 3) begin
					state<=7041;
					out<=115;
				end
				if(in == 4) begin
					state<=3152;
					out<=116;
				end
			end
			5041: begin
				if(in == 0) begin
					state<=5052;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=1154;
					out<=119;
				end
				if(in == 3) begin
					state<=7042;
					out<=120;
				end
				if(in == 4) begin
					state<=3153;
					out<=121;
				end
			end
			5042: begin
				if(in == 0) begin
					state<=5053;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=1155;
					out<=124;
				end
				if(in == 3) begin
					state<=7043;
					out<=125;
				end
				if(in == 4) begin
					state<=3154;
					out<=126;
				end
			end
			5043: begin
				if(in == 0) begin
					state<=5054;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=1156;
					out<=129;
				end
				if(in == 3) begin
					state<=7044;
					out<=130;
				end
				if(in == 4) begin
					state<=3155;
					out<=131;
				end
			end
			5044: begin
				if(in == 0) begin
					state<=5055;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=1157;
					out<=134;
				end
				if(in == 3) begin
					state<=7045;
					out<=135;
				end
				if(in == 4) begin
					state<=3156;
					out<=136;
				end
			end
			5045: begin
				if(in == 0) begin
					state<=5056;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=1158;
					out<=139;
				end
				if(in == 3) begin
					state<=7046;
					out<=140;
				end
				if(in == 4) begin
					state<=3157;
					out<=141;
				end
			end
			5046: begin
				if(in == 0) begin
					state<=5057;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=1159;
					out<=144;
				end
				if(in == 3) begin
					state<=7047;
					out<=145;
				end
				if(in == 4) begin
					state<=3158;
					out<=146;
				end
			end
			5047: begin
				if(in == 0) begin
					state<=5048;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=1150;
					out<=149;
				end
				if(in == 3) begin
					state<=7038;
					out<=150;
				end
				if(in == 4) begin
					state<=3149;
					out<=151;
				end
			end
			5048: begin
				if(in == 0) begin
					state<=5059;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=1161;
					out<=154;
				end
				if(in == 3) begin
					state<=7049;
					out<=155;
				end
				if(in == 4) begin
					state<=3160;
					out<=156;
				end
			end
			5049: begin
				if(in == 0) begin
					state<=5060;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=1162;
					out<=159;
				end
				if(in == 3) begin
					state<=7050;
					out<=160;
				end
				if(in == 4) begin
					state<=3161;
					out<=161;
				end
			end
			5050: begin
				if(in == 0) begin
					state<=5061;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=1163;
					out<=164;
				end
				if(in == 3) begin
					state<=7051;
					out<=165;
				end
				if(in == 4) begin
					state<=3162;
					out<=166;
				end
			end
			5051: begin
				if(in == 0) begin
					state<=5062;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=1164;
					out<=169;
				end
				if(in == 3) begin
					state<=7052;
					out<=170;
				end
				if(in == 4) begin
					state<=3163;
					out<=171;
				end
			end
			5052: begin
				if(in == 0) begin
					state<=5063;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=1165;
					out<=174;
				end
				if(in == 3) begin
					state<=7053;
					out<=175;
				end
				if(in == 4) begin
					state<=3164;
					out<=176;
				end
			end
			5053: begin
				if(in == 0) begin
					state<=5064;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=1166;
					out<=179;
				end
				if(in == 3) begin
					state<=7054;
					out<=180;
				end
				if(in == 4) begin
					state<=3165;
					out<=181;
				end
			end
			5054: begin
				if(in == 0) begin
					state<=5065;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=1167;
					out<=184;
				end
				if(in == 3) begin
					state<=7055;
					out<=185;
				end
				if(in == 4) begin
					state<=3166;
					out<=186;
				end
			end
			5055: begin
				if(in == 0) begin
					state<=5066;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=1168;
					out<=189;
				end
				if(in == 3) begin
					state<=7056;
					out<=190;
				end
				if(in == 4) begin
					state<=3167;
					out<=191;
				end
			end
			5056: begin
				if(in == 0) begin
					state<=5067;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=1169;
					out<=194;
				end
				if(in == 3) begin
					state<=7057;
					out<=195;
				end
				if(in == 4) begin
					state<=3168;
					out<=196;
				end
			end
			5057: begin
				if(in == 0) begin
					state<=5058;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=1160;
					out<=199;
				end
				if(in == 3) begin
					state<=7048;
					out<=200;
				end
				if(in == 4) begin
					state<=3159;
					out<=201;
				end
			end
			5058: begin
				if(in == 0) begin
					state<=5069;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=1171;
					out<=204;
				end
				if(in == 3) begin
					state<=7059;
					out<=205;
				end
				if(in == 4) begin
					state<=3170;
					out<=206;
				end
			end
			5059: begin
				if(in == 0) begin
					state<=5070;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=1172;
					out<=209;
				end
				if(in == 3) begin
					state<=7060;
					out<=210;
				end
				if(in == 4) begin
					state<=3171;
					out<=211;
				end
			end
			5060: begin
				if(in == 0) begin
					state<=5071;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=1173;
					out<=214;
				end
				if(in == 3) begin
					state<=7061;
					out<=215;
				end
				if(in == 4) begin
					state<=3172;
					out<=216;
				end
			end
			5061: begin
				if(in == 0) begin
					state<=5072;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=1174;
					out<=219;
				end
				if(in == 3) begin
					state<=7062;
					out<=220;
				end
				if(in == 4) begin
					state<=3173;
					out<=221;
				end
			end
			5062: begin
				if(in == 0) begin
					state<=5073;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=1175;
					out<=224;
				end
				if(in == 3) begin
					state<=7063;
					out<=225;
				end
				if(in == 4) begin
					state<=3174;
					out<=226;
				end
			end
			5063: begin
				if(in == 0) begin
					state<=5074;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=1176;
					out<=229;
				end
				if(in == 3) begin
					state<=7064;
					out<=230;
				end
				if(in == 4) begin
					state<=3175;
					out<=231;
				end
			end
			5064: begin
				if(in == 0) begin
					state<=5075;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=1177;
					out<=234;
				end
				if(in == 3) begin
					state<=7065;
					out<=235;
				end
				if(in == 4) begin
					state<=3176;
					out<=236;
				end
			end
			5065: begin
				if(in == 0) begin
					state<=5076;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=1178;
					out<=239;
				end
				if(in == 3) begin
					state<=7066;
					out<=240;
				end
				if(in == 4) begin
					state<=3177;
					out<=241;
				end
			end
			5066: begin
				if(in == 0) begin
					state<=5077;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=1179;
					out<=244;
				end
				if(in == 3) begin
					state<=7067;
					out<=245;
				end
				if(in == 4) begin
					state<=3178;
					out<=246;
				end
			end
			5067: begin
				if(in == 0) begin
					state<=5068;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=1170;
					out<=249;
				end
				if(in == 3) begin
					state<=7058;
					out<=250;
				end
				if(in == 4) begin
					state<=3169;
					out<=251;
				end
			end
			5068: begin
				if(in == 0) begin
					state<=5079;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=1181;
					out<=254;
				end
				if(in == 3) begin
					state<=7069;
					out<=255;
				end
				if(in == 4) begin
					state<=3180;
					out<=0;
				end
			end
			5069: begin
				if(in == 0) begin
					state<=5080;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=1182;
					out<=3;
				end
				if(in == 3) begin
					state<=7070;
					out<=4;
				end
				if(in == 4) begin
					state<=3181;
					out<=5;
				end
			end
			5070: begin
				if(in == 0) begin
					state<=5081;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=1183;
					out<=8;
				end
				if(in == 3) begin
					state<=7071;
					out<=9;
				end
				if(in == 4) begin
					state<=3182;
					out<=10;
				end
			end
			5071: begin
				if(in == 0) begin
					state<=5082;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=1184;
					out<=13;
				end
				if(in == 3) begin
					state<=7072;
					out<=14;
				end
				if(in == 4) begin
					state<=3183;
					out<=15;
				end
			end
			5072: begin
				if(in == 0) begin
					state<=5083;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=1185;
					out<=18;
				end
				if(in == 3) begin
					state<=7073;
					out<=19;
				end
				if(in == 4) begin
					state<=3184;
					out<=20;
				end
			end
			5073: begin
				if(in == 0) begin
					state<=5084;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=1186;
					out<=23;
				end
				if(in == 3) begin
					state<=7074;
					out<=24;
				end
				if(in == 4) begin
					state<=3185;
					out<=25;
				end
			end
			5074: begin
				if(in == 0) begin
					state<=5085;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=1187;
					out<=28;
				end
				if(in == 3) begin
					state<=7075;
					out<=29;
				end
				if(in == 4) begin
					state<=3186;
					out<=30;
				end
			end
			5075: begin
				if(in == 0) begin
					state<=5086;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=1188;
					out<=33;
				end
				if(in == 3) begin
					state<=7076;
					out<=34;
				end
				if(in == 4) begin
					state<=3187;
					out<=35;
				end
			end
			5076: begin
				if(in == 0) begin
					state<=5087;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=1189;
					out<=38;
				end
				if(in == 3) begin
					state<=7077;
					out<=39;
				end
				if(in == 4) begin
					state<=3188;
					out<=40;
				end
			end
			5077: begin
				if(in == 0) begin
					state<=5078;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=1180;
					out<=43;
				end
				if(in == 3) begin
					state<=7068;
					out<=44;
				end
				if(in == 4) begin
					state<=3179;
					out<=45;
				end
			end
			5078: begin
				if(in == 0) begin
					state<=5089;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=1191;
					out<=48;
				end
				if(in == 3) begin
					state<=7079;
					out<=49;
				end
				if(in == 4) begin
					state<=3190;
					out<=50;
				end
			end
			5079: begin
				if(in == 0) begin
					state<=5090;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=1192;
					out<=53;
				end
				if(in == 3) begin
					state<=7080;
					out<=54;
				end
				if(in == 4) begin
					state<=3191;
					out<=55;
				end
			end
			5080: begin
				if(in == 0) begin
					state<=5091;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=1193;
					out<=58;
				end
				if(in == 3) begin
					state<=7081;
					out<=59;
				end
				if(in == 4) begin
					state<=3192;
					out<=60;
				end
			end
			5081: begin
				if(in == 0) begin
					state<=5092;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=1194;
					out<=63;
				end
				if(in == 3) begin
					state<=7082;
					out<=64;
				end
				if(in == 4) begin
					state<=3193;
					out<=65;
				end
			end
			5082: begin
				if(in == 0) begin
					state<=5093;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=1195;
					out<=68;
				end
				if(in == 3) begin
					state<=7083;
					out<=69;
				end
				if(in == 4) begin
					state<=3194;
					out<=70;
				end
			end
			5083: begin
				if(in == 0) begin
					state<=5094;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=1196;
					out<=73;
				end
				if(in == 3) begin
					state<=7084;
					out<=74;
				end
				if(in == 4) begin
					state<=3195;
					out<=75;
				end
			end
			5084: begin
				if(in == 0) begin
					state<=5095;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=1197;
					out<=78;
				end
				if(in == 3) begin
					state<=7085;
					out<=79;
				end
				if(in == 4) begin
					state<=3196;
					out<=80;
				end
			end
			5085: begin
				if(in == 0) begin
					state<=5096;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=1198;
					out<=83;
				end
				if(in == 3) begin
					state<=7086;
					out<=84;
				end
				if(in == 4) begin
					state<=3197;
					out<=85;
				end
			end
			5086: begin
				if(in == 0) begin
					state<=5097;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=1199;
					out<=88;
				end
				if(in == 3) begin
					state<=7087;
					out<=89;
				end
				if(in == 4) begin
					state<=3198;
					out<=90;
				end
			end
			5087: begin
				if(in == 0) begin
					state<=5088;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=1190;
					out<=93;
				end
				if(in == 3) begin
					state<=7078;
					out<=94;
				end
				if(in == 4) begin
					state<=3189;
					out<=95;
				end
			end
			5088: begin
				if(in == 0) begin
					state<=5099;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=1201;
					out<=98;
				end
				if(in == 3) begin
					state<=7089;
					out<=99;
				end
				if(in == 4) begin
					state<=3200;
					out<=100;
				end
			end
			5089: begin
				if(in == 0) begin
					state<=5100;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=1202;
					out<=103;
				end
				if(in == 3) begin
					state<=7090;
					out<=104;
				end
				if(in == 4) begin
					state<=3201;
					out<=105;
				end
			end
			5090: begin
				if(in == 0) begin
					state<=5101;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=1203;
					out<=108;
				end
				if(in == 3) begin
					state<=7091;
					out<=109;
				end
				if(in == 4) begin
					state<=3202;
					out<=110;
				end
			end
			5091: begin
				if(in == 0) begin
					state<=5102;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=1204;
					out<=113;
				end
				if(in == 3) begin
					state<=7092;
					out<=114;
				end
				if(in == 4) begin
					state<=3203;
					out<=115;
				end
			end
			5092: begin
				if(in == 0) begin
					state<=5103;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=1205;
					out<=118;
				end
				if(in == 3) begin
					state<=7093;
					out<=119;
				end
				if(in == 4) begin
					state<=3204;
					out<=120;
				end
			end
			5093: begin
				if(in == 0) begin
					state<=5104;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=1206;
					out<=123;
				end
				if(in == 3) begin
					state<=7094;
					out<=124;
				end
				if(in == 4) begin
					state<=3205;
					out<=125;
				end
			end
			5094: begin
				if(in == 0) begin
					state<=5105;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=1207;
					out<=128;
				end
				if(in == 3) begin
					state<=7095;
					out<=129;
				end
				if(in == 4) begin
					state<=3206;
					out<=130;
				end
			end
			5095: begin
				if(in == 0) begin
					state<=5106;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=1208;
					out<=133;
				end
				if(in == 3) begin
					state<=7096;
					out<=134;
				end
				if(in == 4) begin
					state<=3207;
					out<=135;
				end
			end
			5096: begin
				if(in == 0) begin
					state<=5107;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=1209;
					out<=138;
				end
				if(in == 3) begin
					state<=7097;
					out<=139;
				end
				if(in == 4) begin
					state<=3208;
					out<=140;
				end
			end
			5097: begin
				if(in == 0) begin
					state<=5098;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=1200;
					out<=143;
				end
				if(in == 3) begin
					state<=7088;
					out<=144;
				end
				if(in == 4) begin
					state<=3199;
					out<=145;
				end
			end
			5098: begin
				if(in == 0) begin
					state<=5109;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=1211;
					out<=148;
				end
				if(in == 3) begin
					state<=7099;
					out<=149;
				end
				if(in == 4) begin
					state<=3210;
					out<=150;
				end
			end
			5099: begin
				if(in == 0) begin
					state<=5110;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=1212;
					out<=153;
				end
				if(in == 3) begin
					state<=7100;
					out<=154;
				end
				if(in == 4) begin
					state<=3211;
					out<=155;
				end
			end
			5100: begin
				if(in == 0) begin
					state<=5111;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=1213;
					out<=158;
				end
				if(in == 3) begin
					state<=7101;
					out<=159;
				end
				if(in == 4) begin
					state<=3212;
					out<=160;
				end
			end
			5101: begin
				if(in == 0) begin
					state<=5112;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=1214;
					out<=163;
				end
				if(in == 3) begin
					state<=7102;
					out<=164;
				end
				if(in == 4) begin
					state<=3213;
					out<=165;
				end
			end
			5102: begin
				if(in == 0) begin
					state<=5113;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=1215;
					out<=168;
				end
				if(in == 3) begin
					state<=7103;
					out<=169;
				end
				if(in == 4) begin
					state<=3214;
					out<=170;
				end
			end
			5103: begin
				if(in == 0) begin
					state<=5114;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=1216;
					out<=173;
				end
				if(in == 3) begin
					state<=7104;
					out<=174;
				end
				if(in == 4) begin
					state<=3215;
					out<=175;
				end
			end
			5104: begin
				if(in == 0) begin
					state<=5115;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=1217;
					out<=178;
				end
				if(in == 3) begin
					state<=7105;
					out<=179;
				end
				if(in == 4) begin
					state<=3216;
					out<=180;
				end
			end
			5105: begin
				if(in == 0) begin
					state<=5116;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=1218;
					out<=183;
				end
				if(in == 3) begin
					state<=7106;
					out<=184;
				end
				if(in == 4) begin
					state<=3217;
					out<=185;
				end
			end
			5106: begin
				if(in == 0) begin
					state<=5117;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=1219;
					out<=188;
				end
				if(in == 3) begin
					state<=7107;
					out<=189;
				end
				if(in == 4) begin
					state<=3218;
					out<=190;
				end
			end
			5107: begin
				if(in == 0) begin
					state<=5108;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=1210;
					out<=193;
				end
				if(in == 3) begin
					state<=7098;
					out<=194;
				end
				if(in == 4) begin
					state<=3209;
					out<=195;
				end
			end
			5108: begin
				if(in == 0) begin
					state<=5119;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=1221;
					out<=198;
				end
				if(in == 3) begin
					state<=7109;
					out<=199;
				end
				if(in == 4) begin
					state<=3220;
					out<=200;
				end
			end
			5109: begin
				if(in == 0) begin
					state<=5120;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=1222;
					out<=203;
				end
				if(in == 3) begin
					state<=7110;
					out<=204;
				end
				if(in == 4) begin
					state<=3221;
					out<=205;
				end
			end
			5110: begin
				if(in == 0) begin
					state<=5121;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=1223;
					out<=208;
				end
				if(in == 3) begin
					state<=7111;
					out<=209;
				end
				if(in == 4) begin
					state<=3222;
					out<=210;
				end
			end
			5111: begin
				if(in == 0) begin
					state<=5122;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=1224;
					out<=213;
				end
				if(in == 3) begin
					state<=7112;
					out<=214;
				end
				if(in == 4) begin
					state<=3223;
					out<=215;
				end
			end
			5112: begin
				if(in == 0) begin
					state<=5123;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=1225;
					out<=218;
				end
				if(in == 3) begin
					state<=7113;
					out<=219;
				end
				if(in == 4) begin
					state<=3224;
					out<=220;
				end
			end
			5113: begin
				if(in == 0) begin
					state<=5124;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=1226;
					out<=223;
				end
				if(in == 3) begin
					state<=7114;
					out<=224;
				end
				if(in == 4) begin
					state<=3225;
					out<=225;
				end
			end
			5114: begin
				if(in == 0) begin
					state<=5125;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=1227;
					out<=228;
				end
				if(in == 3) begin
					state<=7115;
					out<=229;
				end
				if(in == 4) begin
					state<=3226;
					out<=230;
				end
			end
			5115: begin
				if(in == 0) begin
					state<=5126;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=1228;
					out<=233;
				end
				if(in == 3) begin
					state<=7116;
					out<=234;
				end
				if(in == 4) begin
					state<=3227;
					out<=235;
				end
			end
			5116: begin
				if(in == 0) begin
					state<=5127;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=1229;
					out<=238;
				end
				if(in == 3) begin
					state<=7117;
					out<=239;
				end
				if(in == 4) begin
					state<=3228;
					out<=240;
				end
			end
			5117: begin
				if(in == 0) begin
					state<=5118;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=1220;
					out<=243;
				end
				if(in == 3) begin
					state<=7108;
					out<=244;
				end
				if(in == 4) begin
					state<=3219;
					out<=245;
				end
			end
			5118: begin
				if(in == 0) begin
					state<=4589;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=691;
					out<=248;
				end
				if(in == 3) begin
					state<=6578;
					out<=249;
				end
				if(in == 4) begin
					state<=2689;
					out<=250;
				end
			end
			5119: begin
				if(in == 0) begin
					state<=4590;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=692;
					out<=253;
				end
				if(in == 3) begin
					state<=6579;
					out<=254;
				end
				if(in == 4) begin
					state<=2690;
					out<=255;
				end
			end
			5120: begin
				if(in == 0) begin
					state<=4591;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=693;
					out<=2;
				end
				if(in == 3) begin
					state<=6580;
					out<=3;
				end
				if(in == 4) begin
					state<=2691;
					out<=4;
				end
			end
			5121: begin
				if(in == 0) begin
					state<=4592;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=694;
					out<=7;
				end
				if(in == 3) begin
					state<=6581;
					out<=8;
				end
				if(in == 4) begin
					state<=2692;
					out<=9;
				end
			end
			5122: begin
				if(in == 0) begin
					state<=4593;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=695;
					out<=12;
				end
				if(in == 3) begin
					state<=6582;
					out<=13;
				end
				if(in == 4) begin
					state<=2693;
					out<=14;
				end
			end
			5123: begin
				if(in == 0) begin
					state<=4594;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=696;
					out<=17;
				end
				if(in == 3) begin
					state<=6583;
					out<=18;
				end
				if(in == 4) begin
					state<=2694;
					out<=19;
				end
			end
			5124: begin
				if(in == 0) begin
					state<=4595;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=697;
					out<=22;
				end
				if(in == 3) begin
					state<=6584;
					out<=23;
				end
				if(in == 4) begin
					state<=2695;
					out<=24;
				end
			end
			5125: begin
				if(in == 0) begin
					state<=4596;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=698;
					out<=27;
				end
				if(in == 3) begin
					state<=6585;
					out<=28;
				end
				if(in == 4) begin
					state<=2696;
					out<=29;
				end
			end
			5126: begin
				if(in == 0) begin
					state<=4597;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=699;
					out<=32;
				end
				if(in == 3) begin
					state<=6586;
					out<=33;
				end
				if(in == 4) begin
					state<=2697;
					out<=34;
				end
			end
			5127: begin
				if(in == 0) begin
					state<=5128;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=1230;
					out<=37;
				end
				if(in == 3) begin
					state<=7118;
					out<=38;
				end
				if(in == 4) begin
					state<=3229;
					out<=39;
				end
			end
			5128: begin
				if(in == 0) begin
					state<=4599;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=701;
					out<=42;
				end
				if(in == 3) begin
					state<=6588;
					out<=43;
				end
				if(in == 4) begin
					state<=2699;
					out<=44;
				end
			end
			5129: begin
				if(in == 0) begin
					state<=5140;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=1242;
					out<=47;
				end
				if(in == 3) begin
					state<=6521;
					out<=48;
				end
				if(in == 4) begin
					state<=2632;
					out<=49;
				end
			end
			5130: begin
				if(in == 0) begin
					state<=5141;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=1243;
					out<=52;
				end
				if(in == 3) begin
					state<=6522;
					out<=53;
				end
				if(in == 4) begin
					state<=2633;
					out<=54;
				end
			end
			5131: begin
				if(in == 0) begin
					state<=5142;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=1244;
					out<=57;
				end
				if(in == 3) begin
					state<=6523;
					out<=58;
				end
				if(in == 4) begin
					state<=2634;
					out<=59;
				end
			end
			5132: begin
				if(in == 0) begin
					state<=5143;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=1245;
					out<=62;
				end
				if(in == 3) begin
					state<=6524;
					out<=63;
				end
				if(in == 4) begin
					state<=2635;
					out<=64;
				end
			end
			5133: begin
				if(in == 0) begin
					state<=5144;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=1246;
					out<=67;
				end
				if(in == 3) begin
					state<=6525;
					out<=68;
				end
				if(in == 4) begin
					state<=2636;
					out<=69;
				end
			end
			5134: begin
				if(in == 0) begin
					state<=5145;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=1247;
					out<=72;
				end
				if(in == 3) begin
					state<=6526;
					out<=73;
				end
				if(in == 4) begin
					state<=2637;
					out<=74;
				end
			end
			5135: begin
				if(in == 0) begin
					state<=5146;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=1248;
					out<=77;
				end
				if(in == 3) begin
					state<=6527;
					out<=78;
				end
				if(in == 4) begin
					state<=2638;
					out<=79;
				end
			end
			5136: begin
				if(in == 0) begin
					state<=5147;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=1249;
					out<=82;
				end
				if(in == 3) begin
					state<=6528;
					out<=83;
				end
				if(in == 4) begin
					state<=2639;
					out<=84;
				end
			end
			5137: begin
				if(in == 0) begin
					state<=5138;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=1240;
					out<=87;
				end
				if(in == 3) begin
					state<=6519;
					out<=88;
				end
				if(in == 4) begin
					state<=2630;
					out<=89;
				end
			end
			5138: begin
				if(in == 0) begin
					state<=5149;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=1251;
					out<=92;
				end
				if(in == 3) begin
					state<=6530;
					out<=93;
				end
				if(in == 4) begin
					state<=2641;
					out<=94;
				end
			end
			5139: begin
				if(in == 0) begin
					state<=5150;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=1252;
					out<=97;
				end
				if(in == 3) begin
					state<=6531;
					out<=98;
				end
				if(in == 4) begin
					state<=2642;
					out<=99;
				end
			end
			5140: begin
				if(in == 0) begin
					state<=5151;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=1253;
					out<=102;
				end
				if(in == 3) begin
					state<=6532;
					out<=103;
				end
				if(in == 4) begin
					state<=2643;
					out<=104;
				end
			end
			5141: begin
				if(in == 0) begin
					state<=5152;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=1254;
					out<=107;
				end
				if(in == 3) begin
					state<=6533;
					out<=108;
				end
				if(in == 4) begin
					state<=2644;
					out<=109;
				end
			end
			5142: begin
				if(in == 0) begin
					state<=5153;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=1255;
					out<=112;
				end
				if(in == 3) begin
					state<=6534;
					out<=113;
				end
				if(in == 4) begin
					state<=2645;
					out<=114;
				end
			end
			5143: begin
				if(in == 0) begin
					state<=5154;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=1256;
					out<=117;
				end
				if(in == 3) begin
					state<=6535;
					out<=118;
				end
				if(in == 4) begin
					state<=2646;
					out<=119;
				end
			end
			5144: begin
				if(in == 0) begin
					state<=5155;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=1257;
					out<=122;
				end
				if(in == 3) begin
					state<=6536;
					out<=123;
				end
				if(in == 4) begin
					state<=2647;
					out<=124;
				end
			end
			5145: begin
				if(in == 0) begin
					state<=5156;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=1258;
					out<=127;
				end
				if(in == 3) begin
					state<=6537;
					out<=128;
				end
				if(in == 4) begin
					state<=2648;
					out<=129;
				end
			end
			5146: begin
				if(in == 0) begin
					state<=5157;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=1259;
					out<=132;
				end
				if(in == 3) begin
					state<=6538;
					out<=133;
				end
				if(in == 4) begin
					state<=2649;
					out<=134;
				end
			end
			5147: begin
				if(in == 0) begin
					state<=5148;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=1250;
					out<=137;
				end
				if(in == 3) begin
					state<=6529;
					out<=138;
				end
				if(in == 4) begin
					state<=2640;
					out<=139;
				end
			end
			5148: begin
				if(in == 0) begin
					state<=5159;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=1261;
					out<=142;
				end
				if(in == 3) begin
					state<=6540;
					out<=143;
				end
				if(in == 4) begin
					state<=2651;
					out<=144;
				end
			end
			5149: begin
				if(in == 0) begin
					state<=5160;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=1262;
					out<=147;
				end
				if(in == 3) begin
					state<=6541;
					out<=148;
				end
				if(in == 4) begin
					state<=2652;
					out<=149;
				end
			end
			5150: begin
				if(in == 0) begin
					state<=5161;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=1263;
					out<=152;
				end
				if(in == 3) begin
					state<=6542;
					out<=153;
				end
				if(in == 4) begin
					state<=2653;
					out<=154;
				end
			end
			5151: begin
				if(in == 0) begin
					state<=5162;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=1264;
					out<=157;
				end
				if(in == 3) begin
					state<=6543;
					out<=158;
				end
				if(in == 4) begin
					state<=2654;
					out<=159;
				end
			end
			5152: begin
				if(in == 0) begin
					state<=5163;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=1265;
					out<=162;
				end
				if(in == 3) begin
					state<=6544;
					out<=163;
				end
				if(in == 4) begin
					state<=2655;
					out<=164;
				end
			end
			5153: begin
				if(in == 0) begin
					state<=5164;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=1266;
					out<=167;
				end
				if(in == 3) begin
					state<=6545;
					out<=168;
				end
				if(in == 4) begin
					state<=2656;
					out<=169;
				end
			end
			5154: begin
				if(in == 0) begin
					state<=5165;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=1267;
					out<=172;
				end
				if(in == 3) begin
					state<=6546;
					out<=173;
				end
				if(in == 4) begin
					state<=2657;
					out<=174;
				end
			end
			5155: begin
				if(in == 0) begin
					state<=5166;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=1268;
					out<=177;
				end
				if(in == 3) begin
					state<=6547;
					out<=178;
				end
				if(in == 4) begin
					state<=2658;
					out<=179;
				end
			end
			5156: begin
				if(in == 0) begin
					state<=5167;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=1269;
					out<=182;
				end
				if(in == 3) begin
					state<=6548;
					out<=183;
				end
				if(in == 4) begin
					state<=2659;
					out<=184;
				end
			end
			5157: begin
				if(in == 0) begin
					state<=5158;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=1260;
					out<=187;
				end
				if(in == 3) begin
					state<=6539;
					out<=188;
				end
				if(in == 4) begin
					state<=2650;
					out<=189;
				end
			end
			5158: begin
				if(in == 0) begin
					state<=5169;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=1271;
					out<=192;
				end
				if(in == 3) begin
					state<=6550;
					out<=193;
				end
				if(in == 4) begin
					state<=2661;
					out<=194;
				end
			end
			5159: begin
				if(in == 0) begin
					state<=5170;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=1272;
					out<=197;
				end
				if(in == 3) begin
					state<=6551;
					out<=198;
				end
				if(in == 4) begin
					state<=2662;
					out<=199;
				end
			end
			5160: begin
				if(in == 0) begin
					state<=5171;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=1273;
					out<=202;
				end
				if(in == 3) begin
					state<=6552;
					out<=203;
				end
				if(in == 4) begin
					state<=2663;
					out<=204;
				end
			end
			5161: begin
				if(in == 0) begin
					state<=5172;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=1274;
					out<=207;
				end
				if(in == 3) begin
					state<=6553;
					out<=208;
				end
				if(in == 4) begin
					state<=2664;
					out<=209;
				end
			end
			5162: begin
				if(in == 0) begin
					state<=5173;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=1275;
					out<=212;
				end
				if(in == 3) begin
					state<=6554;
					out<=213;
				end
				if(in == 4) begin
					state<=2665;
					out<=214;
				end
			end
			5163: begin
				if(in == 0) begin
					state<=5174;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=1276;
					out<=217;
				end
				if(in == 3) begin
					state<=6555;
					out<=218;
				end
				if(in == 4) begin
					state<=2666;
					out<=219;
				end
			end
			5164: begin
				if(in == 0) begin
					state<=5175;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=1277;
					out<=222;
				end
				if(in == 3) begin
					state<=6556;
					out<=223;
				end
				if(in == 4) begin
					state<=2667;
					out<=224;
				end
			end
			5165: begin
				if(in == 0) begin
					state<=5176;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=1278;
					out<=227;
				end
				if(in == 3) begin
					state<=6557;
					out<=228;
				end
				if(in == 4) begin
					state<=2668;
					out<=229;
				end
			end
			5166: begin
				if(in == 0) begin
					state<=5177;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=1279;
					out<=232;
				end
				if(in == 3) begin
					state<=6558;
					out<=233;
				end
				if(in == 4) begin
					state<=2669;
					out<=234;
				end
			end
			5167: begin
				if(in == 0) begin
					state<=5168;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=1270;
					out<=237;
				end
				if(in == 3) begin
					state<=6549;
					out<=238;
				end
				if(in == 4) begin
					state<=2660;
					out<=239;
				end
			end
			5168: begin
				if(in == 0) begin
					state<=5179;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=1281;
					out<=242;
				end
				if(in == 3) begin
					state<=7120;
					out<=243;
				end
				if(in == 4) begin
					state<=3231;
					out<=244;
				end
			end
			5169: begin
				if(in == 0) begin
					state<=5180;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=1282;
					out<=247;
				end
				if(in == 3) begin
					state<=7121;
					out<=248;
				end
				if(in == 4) begin
					state<=3232;
					out<=249;
				end
			end
			5170: begin
				if(in == 0) begin
					state<=5181;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=1283;
					out<=252;
				end
				if(in == 3) begin
					state<=7122;
					out<=253;
				end
				if(in == 4) begin
					state<=3233;
					out<=254;
				end
			end
			5171: begin
				if(in == 0) begin
					state<=5182;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=1284;
					out<=1;
				end
				if(in == 3) begin
					state<=7123;
					out<=2;
				end
				if(in == 4) begin
					state<=3234;
					out<=3;
				end
			end
			5172: begin
				if(in == 0) begin
					state<=5183;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=1285;
					out<=6;
				end
				if(in == 3) begin
					state<=7124;
					out<=7;
				end
				if(in == 4) begin
					state<=3235;
					out<=8;
				end
			end
			5173: begin
				if(in == 0) begin
					state<=5184;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=1286;
					out<=11;
				end
				if(in == 3) begin
					state<=7125;
					out<=12;
				end
				if(in == 4) begin
					state<=3236;
					out<=13;
				end
			end
			5174: begin
				if(in == 0) begin
					state<=5185;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=1287;
					out<=16;
				end
				if(in == 3) begin
					state<=7126;
					out<=17;
				end
				if(in == 4) begin
					state<=3237;
					out<=18;
				end
			end
			5175: begin
				if(in == 0) begin
					state<=5186;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=1288;
					out<=21;
				end
				if(in == 3) begin
					state<=7127;
					out<=22;
				end
				if(in == 4) begin
					state<=3238;
					out<=23;
				end
			end
			5176: begin
				if(in == 0) begin
					state<=5187;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=1289;
					out<=26;
				end
				if(in == 3) begin
					state<=7128;
					out<=27;
				end
				if(in == 4) begin
					state<=3239;
					out<=28;
				end
			end
			5177: begin
				if(in == 0) begin
					state<=5178;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=1280;
					out<=31;
				end
				if(in == 3) begin
					state<=7119;
					out<=32;
				end
				if(in == 4) begin
					state<=3230;
					out<=33;
				end
			end
			5178: begin
				if(in == 0) begin
					state<=5189;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=1291;
					out<=36;
				end
				if(in == 3) begin
					state<=7130;
					out<=37;
				end
				if(in == 4) begin
					state<=3241;
					out<=38;
				end
			end
			5179: begin
				if(in == 0) begin
					state<=5190;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=1292;
					out<=41;
				end
				if(in == 3) begin
					state<=7131;
					out<=42;
				end
				if(in == 4) begin
					state<=3242;
					out<=43;
				end
			end
			5180: begin
				if(in == 0) begin
					state<=5191;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=1293;
					out<=46;
				end
				if(in == 3) begin
					state<=7132;
					out<=47;
				end
				if(in == 4) begin
					state<=3243;
					out<=48;
				end
			end
			5181: begin
				if(in == 0) begin
					state<=5192;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=1294;
					out<=51;
				end
				if(in == 3) begin
					state<=7133;
					out<=52;
				end
				if(in == 4) begin
					state<=3244;
					out<=53;
				end
			end
			5182: begin
				if(in == 0) begin
					state<=5193;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=1295;
					out<=56;
				end
				if(in == 3) begin
					state<=7134;
					out<=57;
				end
				if(in == 4) begin
					state<=3245;
					out<=58;
				end
			end
			5183: begin
				if(in == 0) begin
					state<=5194;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=1296;
					out<=61;
				end
				if(in == 3) begin
					state<=7135;
					out<=62;
				end
				if(in == 4) begin
					state<=3246;
					out<=63;
				end
			end
			5184: begin
				if(in == 0) begin
					state<=5195;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=1297;
					out<=66;
				end
				if(in == 3) begin
					state<=7136;
					out<=67;
				end
				if(in == 4) begin
					state<=3247;
					out<=68;
				end
			end
			5185: begin
				if(in == 0) begin
					state<=5196;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=1298;
					out<=71;
				end
				if(in == 3) begin
					state<=7137;
					out<=72;
				end
				if(in == 4) begin
					state<=3248;
					out<=73;
				end
			end
			5186: begin
				if(in == 0) begin
					state<=5197;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=1299;
					out<=76;
				end
				if(in == 3) begin
					state<=7138;
					out<=77;
				end
				if(in == 4) begin
					state<=3249;
					out<=78;
				end
			end
			5187: begin
				if(in == 0) begin
					state<=5188;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=1290;
					out<=81;
				end
				if(in == 3) begin
					state<=7129;
					out<=82;
				end
				if(in == 4) begin
					state<=3240;
					out<=83;
				end
			end
			5188: begin
				if(in == 0) begin
					state<=5199;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=1301;
					out<=86;
				end
				if(in == 3) begin
					state<=7140;
					out<=87;
				end
				if(in == 4) begin
					state<=3251;
					out<=88;
				end
			end
			5189: begin
				if(in == 0) begin
					state<=5200;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=1302;
					out<=91;
				end
				if(in == 3) begin
					state<=7141;
					out<=92;
				end
				if(in == 4) begin
					state<=3252;
					out<=93;
				end
			end
			5190: begin
				if(in == 0) begin
					state<=5201;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=1303;
					out<=96;
				end
				if(in == 3) begin
					state<=7142;
					out<=97;
				end
				if(in == 4) begin
					state<=3253;
					out<=98;
				end
			end
			5191: begin
				if(in == 0) begin
					state<=5202;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=1304;
					out<=101;
				end
				if(in == 3) begin
					state<=7143;
					out<=102;
				end
				if(in == 4) begin
					state<=3254;
					out<=103;
				end
			end
			5192: begin
				if(in == 0) begin
					state<=5203;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=1305;
					out<=106;
				end
				if(in == 3) begin
					state<=7144;
					out<=107;
				end
				if(in == 4) begin
					state<=3255;
					out<=108;
				end
			end
			5193: begin
				if(in == 0) begin
					state<=5204;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=1306;
					out<=111;
				end
				if(in == 3) begin
					state<=7145;
					out<=112;
				end
				if(in == 4) begin
					state<=3256;
					out<=113;
				end
			end
			5194: begin
				if(in == 0) begin
					state<=5205;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=1307;
					out<=116;
				end
				if(in == 3) begin
					state<=7146;
					out<=117;
				end
				if(in == 4) begin
					state<=3257;
					out<=118;
				end
			end
			5195: begin
				if(in == 0) begin
					state<=5206;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=1308;
					out<=121;
				end
				if(in == 3) begin
					state<=7147;
					out<=122;
				end
				if(in == 4) begin
					state<=3258;
					out<=123;
				end
			end
			5196: begin
				if(in == 0) begin
					state<=5207;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=1309;
					out<=126;
				end
				if(in == 3) begin
					state<=7148;
					out<=127;
				end
				if(in == 4) begin
					state<=3259;
					out<=128;
				end
			end
			5197: begin
				if(in == 0) begin
					state<=5198;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=1300;
					out<=131;
				end
				if(in == 3) begin
					state<=7139;
					out<=132;
				end
				if(in == 4) begin
					state<=3250;
					out<=133;
				end
			end
			5198: begin
				if(in == 0) begin
					state<=5209;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=1311;
					out<=136;
				end
				if(in == 3) begin
					state<=6559;
					out<=137;
				end
				if(in == 4) begin
					state<=2670;
					out<=138;
				end
			end
			5199: begin
				if(in == 0) begin
					state<=5210;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=1312;
					out<=141;
				end
				if(in == 3) begin
					state<=6560;
					out<=142;
				end
				if(in == 4) begin
					state<=2671;
					out<=143;
				end
			end
			5200: begin
				if(in == 0) begin
					state<=5211;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=1313;
					out<=146;
				end
				if(in == 3) begin
					state<=6561;
					out<=147;
				end
				if(in == 4) begin
					state<=2672;
					out<=148;
				end
			end
			5201: begin
				if(in == 0) begin
					state<=5212;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=1314;
					out<=151;
				end
				if(in == 3) begin
					state<=6562;
					out<=152;
				end
				if(in == 4) begin
					state<=2673;
					out<=153;
				end
			end
			5202: begin
				if(in == 0) begin
					state<=5213;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=1315;
					out<=156;
				end
				if(in == 3) begin
					state<=6563;
					out<=157;
				end
				if(in == 4) begin
					state<=2674;
					out<=158;
				end
			end
			5203: begin
				if(in == 0) begin
					state<=5214;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=1316;
					out<=161;
				end
				if(in == 3) begin
					state<=6564;
					out<=162;
				end
				if(in == 4) begin
					state<=2675;
					out<=163;
				end
			end
			5204: begin
				if(in == 0) begin
					state<=5215;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=1317;
					out<=166;
				end
				if(in == 3) begin
					state<=6565;
					out<=167;
				end
				if(in == 4) begin
					state<=2676;
					out<=168;
				end
			end
			5205: begin
				if(in == 0) begin
					state<=5216;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=1318;
					out<=171;
				end
				if(in == 3) begin
					state<=6566;
					out<=172;
				end
				if(in == 4) begin
					state<=2677;
					out<=173;
				end
			end
			5206: begin
				if(in == 0) begin
					state<=5217;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=1319;
					out<=176;
				end
				if(in == 3) begin
					state<=6567;
					out<=177;
				end
				if(in == 4) begin
					state<=2678;
					out<=178;
				end
			end
			5207: begin
				if(in == 0) begin
					state<=5208;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=1310;
					out<=181;
				end
				if(in == 3) begin
					state<=7149;
					out<=182;
				end
				if(in == 4) begin
					state<=3260;
					out<=183;
				end
			end
			5208: begin
				if(in == 0) begin
					state<=4789;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=1321;
					out<=186;
				end
				if(in == 3) begin
					state<=6569;
					out<=187;
				end
				if(in == 4) begin
					state<=2680;
					out<=188;
				end
			end
			5209: begin
				if(in == 0) begin
					state<=4790;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=1322;
					out<=191;
				end
				if(in == 3) begin
					state<=6570;
					out<=192;
				end
				if(in == 4) begin
					state<=2681;
					out<=193;
				end
			end
			5210: begin
				if(in == 0) begin
					state<=4791;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=1323;
					out<=196;
				end
				if(in == 3) begin
					state<=6571;
					out<=197;
				end
				if(in == 4) begin
					state<=2682;
					out<=198;
				end
			end
			5211: begin
				if(in == 0) begin
					state<=4792;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=1324;
					out<=201;
				end
				if(in == 3) begin
					state<=6572;
					out<=202;
				end
				if(in == 4) begin
					state<=2683;
					out<=203;
				end
			end
			5212: begin
				if(in == 0) begin
					state<=4793;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=1325;
					out<=206;
				end
				if(in == 3) begin
					state<=6573;
					out<=207;
				end
				if(in == 4) begin
					state<=2684;
					out<=208;
				end
			end
			5213: begin
				if(in == 0) begin
					state<=4794;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=1326;
					out<=211;
				end
				if(in == 3) begin
					state<=6574;
					out<=212;
				end
				if(in == 4) begin
					state<=2685;
					out<=213;
				end
			end
			5214: begin
				if(in == 0) begin
					state<=4795;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=1327;
					out<=216;
				end
				if(in == 3) begin
					state<=6575;
					out<=217;
				end
				if(in == 4) begin
					state<=2686;
					out<=218;
				end
			end
			5215: begin
				if(in == 0) begin
					state<=4796;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=1328;
					out<=221;
				end
				if(in == 3) begin
					state<=6576;
					out<=222;
				end
				if(in == 4) begin
					state<=2687;
					out<=223;
				end
			end
			5216: begin
				if(in == 0) begin
					state<=4797;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=899;
					out<=226;
				end
				if(in == 3) begin
					state<=6577;
					out<=227;
				end
				if(in == 4) begin
					state<=2688;
					out<=228;
				end
			end
			5217: begin
				if(in == 0) begin
					state<=4788;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=1320;
					out<=231;
				end
				if(in == 3) begin
					state<=6568;
					out<=232;
				end
				if(in == 4) begin
					state<=2679;
					out<=233;
				end
			end
			5218: begin
				if(in == 0) begin
					state<=5229;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=1340;
					out<=236;
				end
				if(in == 3) begin
					state<=7161;
					out<=237;
				end
				if(in == 4) begin
					state<=3272;
					out<=238;
				end
			end
			5219: begin
				if(in == 0) begin
					state<=5230;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=1341;
					out<=241;
				end
				if(in == 3) begin
					state<=7162;
					out<=242;
				end
				if(in == 4) begin
					state<=3273;
					out<=243;
				end
			end
			5220: begin
				if(in == 0) begin
					state<=5231;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=1342;
					out<=246;
				end
				if(in == 3) begin
					state<=7163;
					out<=247;
				end
				if(in == 4) begin
					state<=3274;
					out<=248;
				end
			end
			5221: begin
				if(in == 0) begin
					state<=5232;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=1343;
					out<=251;
				end
				if(in == 3) begin
					state<=7164;
					out<=252;
				end
				if(in == 4) begin
					state<=3275;
					out<=253;
				end
			end
			5222: begin
				if(in == 0) begin
					state<=5233;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=1344;
					out<=0;
				end
				if(in == 3) begin
					state<=7165;
					out<=1;
				end
				if(in == 4) begin
					state<=3276;
					out<=2;
				end
			end
			5223: begin
				if(in == 0) begin
					state<=5234;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=1345;
					out<=5;
				end
				if(in == 3) begin
					state<=7166;
					out<=6;
				end
				if(in == 4) begin
					state<=3277;
					out<=7;
				end
			end
			5224: begin
				if(in == 0) begin
					state<=5235;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=1346;
					out<=10;
				end
				if(in == 3) begin
					state<=7167;
					out<=11;
				end
				if(in == 4) begin
					state<=3278;
					out<=12;
				end
			end
			5225: begin
				if(in == 0) begin
					state<=5236;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=1347;
					out<=15;
				end
				if(in == 3) begin
					state<=7168;
					out<=16;
				end
				if(in == 4) begin
					state<=3279;
					out<=17;
				end
			end
			5226: begin
				if(in == 0) begin
					state<=5237;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=1348;
					out<=20;
				end
				if(in == 3) begin
					state<=7169;
					out<=21;
				end
				if(in == 4) begin
					state<=3280;
					out<=22;
				end
			end
			5227: begin
				if(in == 0) begin
					state<=5228;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=1339;
					out<=25;
				end
				if(in == 3) begin
					state<=7160;
					out<=26;
				end
				if(in == 4) begin
					state<=3271;
					out<=27;
				end
			end
			5228: begin
				if(in == 0) begin
					state<=5239;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=1350;
					out<=30;
				end
				if(in == 3) begin
					state<=7171;
					out<=31;
				end
				if(in == 4) begin
					state<=3282;
					out<=32;
				end
			end
			5229: begin
				if(in == 0) begin
					state<=5240;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=1351;
					out<=35;
				end
				if(in == 3) begin
					state<=7172;
					out<=36;
				end
				if(in == 4) begin
					state<=3283;
					out<=37;
				end
			end
			5230: begin
				if(in == 0) begin
					state<=5241;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=1352;
					out<=40;
				end
				if(in == 3) begin
					state<=7173;
					out<=41;
				end
				if(in == 4) begin
					state<=3284;
					out<=42;
				end
			end
			5231: begin
				if(in == 0) begin
					state<=5242;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=1353;
					out<=45;
				end
				if(in == 3) begin
					state<=7174;
					out<=46;
				end
				if(in == 4) begin
					state<=3285;
					out<=47;
				end
			end
			5232: begin
				if(in == 0) begin
					state<=5243;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=1354;
					out<=50;
				end
				if(in == 3) begin
					state<=7175;
					out<=51;
				end
				if(in == 4) begin
					state<=3286;
					out<=52;
				end
			end
			5233: begin
				if(in == 0) begin
					state<=5244;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=1355;
					out<=55;
				end
				if(in == 3) begin
					state<=7176;
					out<=56;
				end
				if(in == 4) begin
					state<=3287;
					out<=57;
				end
			end
			5234: begin
				if(in == 0) begin
					state<=5245;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=1356;
					out<=60;
				end
				if(in == 3) begin
					state<=7177;
					out<=61;
				end
				if(in == 4) begin
					state<=3288;
					out<=62;
				end
			end
			5235: begin
				if(in == 0) begin
					state<=5246;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=1357;
					out<=65;
				end
				if(in == 3) begin
					state<=7178;
					out<=66;
				end
				if(in == 4) begin
					state<=3289;
					out<=67;
				end
			end
			5236: begin
				if(in == 0) begin
					state<=5247;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=1358;
					out<=70;
				end
				if(in == 3) begin
					state<=7179;
					out<=71;
				end
				if(in == 4) begin
					state<=3290;
					out<=72;
				end
			end
			5237: begin
				if(in == 0) begin
					state<=5238;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=1349;
					out<=75;
				end
				if(in == 3) begin
					state<=7170;
					out<=76;
				end
				if(in == 4) begin
					state<=3281;
					out<=77;
				end
			end
			5238: begin
				if(in == 0) begin
					state<=3949;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=51;
					out<=80;
				end
				if(in == 3) begin
					state<=5938;
					out<=81;
				end
				if(in == 4) begin
					state<=2049;
					out<=82;
				end
			end
			5239: begin
				if(in == 0) begin
					state<=3950;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=52;
					out<=85;
				end
				if(in == 3) begin
					state<=5939;
					out<=86;
				end
				if(in == 4) begin
					state<=2050;
					out<=87;
				end
			end
			5240: begin
				if(in == 0) begin
					state<=3951;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=53;
					out<=90;
				end
				if(in == 3) begin
					state<=5940;
					out<=91;
				end
				if(in == 4) begin
					state<=2051;
					out<=92;
				end
			end
			5241: begin
				if(in == 0) begin
					state<=3952;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=54;
					out<=95;
				end
				if(in == 3) begin
					state<=5941;
					out<=96;
				end
				if(in == 4) begin
					state<=2052;
					out<=97;
				end
			end
			5242: begin
				if(in == 0) begin
					state<=3953;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=55;
					out<=100;
				end
				if(in == 3) begin
					state<=5942;
					out<=101;
				end
				if(in == 4) begin
					state<=2053;
					out<=102;
				end
			end
			5243: begin
				if(in == 0) begin
					state<=3954;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=56;
					out<=105;
				end
				if(in == 3) begin
					state<=5943;
					out<=106;
				end
				if(in == 4) begin
					state<=2054;
					out<=107;
				end
			end
			5244: begin
				if(in == 0) begin
					state<=3955;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=57;
					out<=110;
				end
				if(in == 3) begin
					state<=5944;
					out<=111;
				end
				if(in == 4) begin
					state<=2055;
					out<=112;
				end
			end
			5245: begin
				if(in == 0) begin
					state<=3956;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=58;
					out<=115;
				end
				if(in == 3) begin
					state<=5945;
					out<=116;
				end
				if(in == 4) begin
					state<=2056;
					out<=117;
				end
			end
			5246: begin
				if(in == 0) begin
					state<=3957;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=59;
					out<=120;
				end
				if(in == 3) begin
					state<=5946;
					out<=121;
				end
				if(in == 4) begin
					state<=2057;
					out<=122;
				end
			end
			5247: begin
				if(in == 0) begin
					state<=5248;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=1359;
					out<=125;
				end
				if(in == 3) begin
					state<=7180;
					out<=126;
				end
				if(in == 4) begin
					state<=3291;
					out<=127;
				end
			end
			5248: begin
				if(in == 0) begin
					state<=3959;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=61;
					out<=130;
				end
				if(in == 3) begin
					state<=5948;
					out<=131;
				end
				if(in == 4) begin
					state<=2059;
					out<=132;
				end
			end
			5249: begin
				if(in == 0) begin
					state<=5260;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=1371;
					out<=135;
				end
				if(in == 3) begin
					state<=7192;
					out<=136;
				end
				if(in == 4) begin
					state<=3303;
					out<=137;
				end
			end
			5250: begin
				if(in == 0) begin
					state<=5261;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=1372;
					out<=140;
				end
				if(in == 3) begin
					state<=7193;
					out<=141;
				end
				if(in == 4) begin
					state<=3304;
					out<=142;
				end
			end
			5251: begin
				if(in == 0) begin
					state<=5262;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=1373;
					out<=145;
				end
				if(in == 3) begin
					state<=7194;
					out<=146;
				end
				if(in == 4) begin
					state<=3305;
					out<=147;
				end
			end
			5252: begin
				if(in == 0) begin
					state<=5263;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=1374;
					out<=150;
				end
				if(in == 3) begin
					state<=7195;
					out<=151;
				end
				if(in == 4) begin
					state<=3306;
					out<=152;
				end
			end
			5253: begin
				if(in == 0) begin
					state<=5264;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=1375;
					out<=155;
				end
				if(in == 3) begin
					state<=7196;
					out<=156;
				end
				if(in == 4) begin
					state<=3307;
					out<=157;
				end
			end
			5254: begin
				if(in == 0) begin
					state<=5265;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=1376;
					out<=160;
				end
				if(in == 3) begin
					state<=7197;
					out<=161;
				end
				if(in == 4) begin
					state<=3308;
					out<=162;
				end
			end
			5255: begin
				if(in == 0) begin
					state<=5266;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=1377;
					out<=165;
				end
				if(in == 3) begin
					state<=7198;
					out<=166;
				end
				if(in == 4) begin
					state<=3309;
					out<=167;
				end
			end
			5256: begin
				if(in == 0) begin
					state<=5267;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=1378;
					out<=170;
				end
				if(in == 3) begin
					state<=7199;
					out<=171;
				end
				if(in == 4) begin
					state<=3310;
					out<=172;
				end
			end
			5257: begin
				if(in == 0) begin
					state<=5268;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=1379;
					out<=175;
				end
				if(in == 3) begin
					state<=7200;
					out<=176;
				end
				if(in == 4) begin
					state<=3311;
					out<=177;
				end
			end
			5258: begin
				if(in == 0) begin
					state<=5259;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=1370;
					out<=180;
				end
				if(in == 3) begin
					state<=7191;
					out<=181;
				end
				if(in == 4) begin
					state<=3302;
					out<=182;
				end
			end
			5259: begin
				if(in == 0) begin
					state<=5270;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=1381;
					out<=185;
				end
				if(in == 3) begin
					state<=7202;
					out<=186;
				end
				if(in == 4) begin
					state<=3313;
					out<=187;
				end
			end
			5260: begin
				if(in == 0) begin
					state<=5271;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=1382;
					out<=190;
				end
				if(in == 3) begin
					state<=7203;
					out<=191;
				end
				if(in == 4) begin
					state<=3314;
					out<=192;
				end
			end
			5261: begin
				if(in == 0) begin
					state<=5272;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=1383;
					out<=195;
				end
				if(in == 3) begin
					state<=7204;
					out<=196;
				end
				if(in == 4) begin
					state<=3315;
					out<=197;
				end
			end
			5262: begin
				if(in == 0) begin
					state<=5273;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=1384;
					out<=200;
				end
				if(in == 3) begin
					state<=7205;
					out<=201;
				end
				if(in == 4) begin
					state<=3316;
					out<=202;
				end
			end
			5263: begin
				if(in == 0) begin
					state<=5274;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=1385;
					out<=205;
				end
				if(in == 3) begin
					state<=7206;
					out<=206;
				end
				if(in == 4) begin
					state<=3317;
					out<=207;
				end
			end
			5264: begin
				if(in == 0) begin
					state<=5275;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=1386;
					out<=210;
				end
				if(in == 3) begin
					state<=7207;
					out<=211;
				end
				if(in == 4) begin
					state<=3318;
					out<=212;
				end
			end
			5265: begin
				if(in == 0) begin
					state<=5276;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=1387;
					out<=215;
				end
				if(in == 3) begin
					state<=7208;
					out<=216;
				end
				if(in == 4) begin
					state<=3319;
					out<=217;
				end
			end
			5266: begin
				if(in == 0) begin
					state<=5277;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=1388;
					out<=220;
				end
				if(in == 3) begin
					state<=7209;
					out<=221;
				end
				if(in == 4) begin
					state<=3320;
					out<=222;
				end
			end
			5267: begin
				if(in == 0) begin
					state<=5278;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=1389;
					out<=225;
				end
				if(in == 3) begin
					state<=7210;
					out<=226;
				end
				if(in == 4) begin
					state<=3321;
					out<=227;
				end
			end
			5268: begin
				if(in == 0) begin
					state<=5269;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=1380;
					out<=230;
				end
				if(in == 3) begin
					state<=7201;
					out<=231;
				end
				if(in == 4) begin
					state<=3312;
					out<=232;
				end
			end
			5269: begin
				if(in == 0) begin
					state<=4018;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=120;
					out<=235;
				end
				if(in == 3) begin
					state<=6007;
					out<=236;
				end
				if(in == 4) begin
					state<=2118;
					out<=237;
				end
			end
			5270: begin
				if(in == 0) begin
					state<=4019;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=121;
					out<=240;
				end
				if(in == 3) begin
					state<=6008;
					out<=241;
				end
				if(in == 4) begin
					state<=2119;
					out<=242;
				end
			end
			5271: begin
				if(in == 0) begin
					state<=4020;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=122;
					out<=245;
				end
				if(in == 3) begin
					state<=6009;
					out<=246;
				end
				if(in == 4) begin
					state<=2120;
					out<=247;
				end
			end
			5272: begin
				if(in == 0) begin
					state<=4021;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=123;
					out<=250;
				end
				if(in == 3) begin
					state<=6010;
					out<=251;
				end
				if(in == 4) begin
					state<=2121;
					out<=252;
				end
			end
			5273: begin
				if(in == 0) begin
					state<=4022;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=124;
					out<=255;
				end
				if(in == 3) begin
					state<=6011;
					out<=0;
				end
				if(in == 4) begin
					state<=2122;
					out<=1;
				end
			end
			5274: begin
				if(in == 0) begin
					state<=4023;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=125;
					out<=4;
				end
				if(in == 3) begin
					state<=6012;
					out<=5;
				end
				if(in == 4) begin
					state<=2123;
					out<=6;
				end
			end
			5275: begin
				if(in == 0) begin
					state<=4024;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=126;
					out<=9;
				end
				if(in == 3) begin
					state<=6013;
					out<=10;
				end
				if(in == 4) begin
					state<=2124;
					out<=11;
				end
			end
			5276: begin
				if(in == 0) begin
					state<=4025;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=127;
					out<=14;
				end
				if(in == 3) begin
					state<=6014;
					out<=15;
				end
				if(in == 4) begin
					state<=2125;
					out<=16;
				end
			end
			5277: begin
				if(in == 0) begin
					state<=4026;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=128;
					out<=19;
				end
				if(in == 3) begin
					state<=6015;
					out<=20;
				end
				if(in == 4) begin
					state<=2126;
					out<=21;
				end
			end
			5278: begin
				if(in == 0) begin
					state<=5279;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=1390;
					out<=24;
				end
				if(in == 3) begin
					state<=7211;
					out<=25;
				end
				if(in == 4) begin
					state<=3322;
					out<=26;
				end
			end
			5279: begin
				if(in == 0) begin
					state<=4028;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=130;
					out<=29;
				end
				if(in == 3) begin
					state<=6017;
					out<=30;
				end
				if(in == 4) begin
					state<=2128;
					out<=31;
				end
			end
			5280: begin
				if(in == 0) begin
					state<=5291;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=1402;
					out<=34;
				end
				if(in == 3) begin
					state<=7223;
					out<=35;
				end
				if(in == 4) begin
					state<=3334;
					out<=36;
				end
			end
			5281: begin
				if(in == 0) begin
					state<=5292;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=1403;
					out<=39;
				end
				if(in == 3) begin
					state<=7224;
					out<=40;
				end
				if(in == 4) begin
					state<=3335;
					out<=41;
				end
			end
			5282: begin
				if(in == 0) begin
					state<=5293;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=1404;
					out<=44;
				end
				if(in == 3) begin
					state<=7225;
					out<=45;
				end
				if(in == 4) begin
					state<=3336;
					out<=46;
				end
			end
			5283: begin
				if(in == 0) begin
					state<=5294;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=1405;
					out<=49;
				end
				if(in == 3) begin
					state<=7226;
					out<=50;
				end
				if(in == 4) begin
					state<=3337;
					out<=51;
				end
			end
			5284: begin
				if(in == 0) begin
					state<=5295;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=1406;
					out<=54;
				end
				if(in == 3) begin
					state<=7227;
					out<=55;
				end
				if(in == 4) begin
					state<=3338;
					out<=56;
				end
			end
			5285: begin
				if(in == 0) begin
					state<=5296;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=1407;
					out<=59;
				end
				if(in == 3) begin
					state<=7228;
					out<=60;
				end
				if(in == 4) begin
					state<=3339;
					out<=61;
				end
			end
			5286: begin
				if(in == 0) begin
					state<=5297;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=1408;
					out<=64;
				end
				if(in == 3) begin
					state<=7229;
					out<=65;
				end
				if(in == 4) begin
					state<=3340;
					out<=66;
				end
			end
			5287: begin
				if(in == 0) begin
					state<=5298;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=1409;
					out<=69;
				end
				if(in == 3) begin
					state<=7230;
					out<=70;
				end
				if(in == 4) begin
					state<=3341;
					out<=71;
				end
			end
			5288: begin
				if(in == 0) begin
					state<=5299;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=1410;
					out<=74;
				end
				if(in == 3) begin
					state<=7231;
					out<=75;
				end
				if(in == 4) begin
					state<=3342;
					out<=76;
				end
			end
			5289: begin
				if(in == 0) begin
					state<=5290;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=1401;
					out<=79;
				end
				if(in == 3) begin
					state<=7222;
					out<=80;
				end
				if(in == 4) begin
					state<=3333;
					out<=81;
				end
			end
			5290: begin
				if(in == 0) begin
					state<=5301;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=1412;
					out<=84;
				end
				if(in == 3) begin
					state<=7233;
					out<=85;
				end
				if(in == 4) begin
					state<=3344;
					out<=86;
				end
			end
			5291: begin
				if(in == 0) begin
					state<=5302;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=1413;
					out<=89;
				end
				if(in == 3) begin
					state<=7234;
					out<=90;
				end
				if(in == 4) begin
					state<=3345;
					out<=91;
				end
			end
			5292: begin
				if(in == 0) begin
					state<=5303;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=1414;
					out<=94;
				end
				if(in == 3) begin
					state<=7235;
					out<=95;
				end
				if(in == 4) begin
					state<=3346;
					out<=96;
				end
			end
			5293: begin
				if(in == 0) begin
					state<=5304;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=1415;
					out<=99;
				end
				if(in == 3) begin
					state<=7236;
					out<=100;
				end
				if(in == 4) begin
					state<=3347;
					out<=101;
				end
			end
			5294: begin
				if(in == 0) begin
					state<=5305;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=1416;
					out<=104;
				end
				if(in == 3) begin
					state<=7237;
					out<=105;
				end
				if(in == 4) begin
					state<=3348;
					out<=106;
				end
			end
			5295: begin
				if(in == 0) begin
					state<=5306;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=1417;
					out<=109;
				end
				if(in == 3) begin
					state<=7238;
					out<=110;
				end
				if(in == 4) begin
					state<=3349;
					out<=111;
				end
			end
			5296: begin
				if(in == 0) begin
					state<=5307;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=1418;
					out<=114;
				end
				if(in == 3) begin
					state<=7239;
					out<=115;
				end
				if(in == 4) begin
					state<=3350;
					out<=116;
				end
			end
			5297: begin
				if(in == 0) begin
					state<=5308;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=1419;
					out<=119;
				end
				if(in == 3) begin
					state<=7240;
					out<=120;
				end
				if(in == 4) begin
					state<=3351;
					out<=121;
				end
			end
			5298: begin
				if(in == 0) begin
					state<=5309;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=1420;
					out<=124;
				end
				if(in == 3) begin
					state<=7241;
					out<=125;
				end
				if(in == 4) begin
					state<=3352;
					out<=126;
				end
			end
			5299: begin
				if(in == 0) begin
					state<=5300;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=1411;
					out<=129;
				end
				if(in == 3) begin
					state<=7232;
					out<=130;
				end
				if(in == 4) begin
					state<=3343;
					out<=131;
				end
			end
			5300: begin
				if(in == 0) begin
					state<=4087;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=189;
					out<=134;
				end
				if(in == 3) begin
					state<=6076;
					out<=135;
				end
				if(in == 4) begin
					state<=2187;
					out<=136;
				end
			end
			5301: begin
				if(in == 0) begin
					state<=4088;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=190;
					out<=139;
				end
				if(in == 3) begin
					state<=6077;
					out<=140;
				end
				if(in == 4) begin
					state<=2188;
					out<=141;
				end
			end
			5302: begin
				if(in == 0) begin
					state<=4089;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=191;
					out<=144;
				end
				if(in == 3) begin
					state<=6078;
					out<=145;
				end
				if(in == 4) begin
					state<=2189;
					out<=146;
				end
			end
			5303: begin
				if(in == 0) begin
					state<=4090;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=192;
					out<=149;
				end
				if(in == 3) begin
					state<=6079;
					out<=150;
				end
				if(in == 4) begin
					state<=2190;
					out<=151;
				end
			end
			5304: begin
				if(in == 0) begin
					state<=4091;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=193;
					out<=154;
				end
				if(in == 3) begin
					state<=6080;
					out<=155;
				end
				if(in == 4) begin
					state<=2191;
					out<=156;
				end
			end
			5305: begin
				if(in == 0) begin
					state<=4092;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=194;
					out<=159;
				end
				if(in == 3) begin
					state<=6081;
					out<=160;
				end
				if(in == 4) begin
					state<=2192;
					out<=161;
				end
			end
			5306: begin
				if(in == 0) begin
					state<=4093;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=195;
					out<=164;
				end
				if(in == 3) begin
					state<=6082;
					out<=165;
				end
				if(in == 4) begin
					state<=2193;
					out<=166;
				end
			end
			5307: begin
				if(in == 0) begin
					state<=4094;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=196;
					out<=169;
				end
				if(in == 3) begin
					state<=6083;
					out<=170;
				end
				if(in == 4) begin
					state<=2194;
					out<=171;
				end
			end
			5308: begin
				if(in == 0) begin
					state<=4095;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=197;
					out<=174;
				end
				if(in == 3) begin
					state<=6084;
					out<=175;
				end
				if(in == 4) begin
					state<=2195;
					out<=176;
				end
			end
			5309: begin
				if(in == 0) begin
					state<=5310;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=1421;
					out<=179;
				end
				if(in == 3) begin
					state<=7242;
					out<=180;
				end
				if(in == 4) begin
					state<=3353;
					out<=181;
				end
			end
			5310: begin
				if(in == 0) begin
					state<=4097;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=199;
					out<=184;
				end
				if(in == 3) begin
					state<=6086;
					out<=185;
				end
				if(in == 4) begin
					state<=2197;
					out<=186;
				end
			end
			5311: begin
				if(in == 0) begin
					state<=5322;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=1433;
					out<=189;
				end
				if(in == 3) begin
					state<=7254;
					out<=190;
				end
				if(in == 4) begin
					state<=3365;
					out<=191;
				end
			end
			5312: begin
				if(in == 0) begin
					state<=5323;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=1434;
					out<=194;
				end
				if(in == 3) begin
					state<=7255;
					out<=195;
				end
				if(in == 4) begin
					state<=3366;
					out<=196;
				end
			end
			5313: begin
				if(in == 0) begin
					state<=5324;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=1435;
					out<=199;
				end
				if(in == 3) begin
					state<=7256;
					out<=200;
				end
				if(in == 4) begin
					state<=3367;
					out<=201;
				end
			end
			5314: begin
				if(in == 0) begin
					state<=5325;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=1436;
					out<=204;
				end
				if(in == 3) begin
					state<=7257;
					out<=205;
				end
				if(in == 4) begin
					state<=3368;
					out<=206;
				end
			end
			5315: begin
				if(in == 0) begin
					state<=5326;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=1437;
					out<=209;
				end
				if(in == 3) begin
					state<=7258;
					out<=210;
				end
				if(in == 4) begin
					state<=3369;
					out<=211;
				end
			end
			5316: begin
				if(in == 0) begin
					state<=5327;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=1438;
					out<=214;
				end
				if(in == 3) begin
					state<=7259;
					out<=215;
				end
				if(in == 4) begin
					state<=3370;
					out<=216;
				end
			end
			5317: begin
				if(in == 0) begin
					state<=5328;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=1439;
					out<=219;
				end
				if(in == 3) begin
					state<=7260;
					out<=220;
				end
				if(in == 4) begin
					state<=3371;
					out<=221;
				end
			end
			5318: begin
				if(in == 0) begin
					state<=5329;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=1440;
					out<=224;
				end
				if(in == 3) begin
					state<=7261;
					out<=225;
				end
				if(in == 4) begin
					state<=3372;
					out<=226;
				end
			end
			5319: begin
				if(in == 0) begin
					state<=5330;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=1441;
					out<=229;
				end
				if(in == 3) begin
					state<=7262;
					out<=230;
				end
				if(in == 4) begin
					state<=3373;
					out<=231;
				end
			end
			5320: begin
				if(in == 0) begin
					state<=5321;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=1432;
					out<=234;
				end
				if(in == 3) begin
					state<=7253;
					out<=235;
				end
				if(in == 4) begin
					state<=3364;
					out<=236;
				end
			end
			5321: begin
				if(in == 0) begin
					state<=5332;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=1443;
					out<=239;
				end
				if(in == 3) begin
					state<=7264;
					out<=240;
				end
				if(in == 4) begin
					state<=3375;
					out<=241;
				end
			end
			5322: begin
				if(in == 0) begin
					state<=5333;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=1444;
					out<=244;
				end
				if(in == 3) begin
					state<=7265;
					out<=245;
				end
				if(in == 4) begin
					state<=3376;
					out<=246;
				end
			end
			5323: begin
				if(in == 0) begin
					state<=5334;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=1445;
					out<=249;
				end
				if(in == 3) begin
					state<=7266;
					out<=250;
				end
				if(in == 4) begin
					state<=3377;
					out<=251;
				end
			end
			5324: begin
				if(in == 0) begin
					state<=5335;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=1446;
					out<=254;
				end
				if(in == 3) begin
					state<=7267;
					out<=255;
				end
				if(in == 4) begin
					state<=3378;
					out<=0;
				end
			end
			5325: begin
				if(in == 0) begin
					state<=5336;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=1447;
					out<=3;
				end
				if(in == 3) begin
					state<=7268;
					out<=4;
				end
				if(in == 4) begin
					state<=3379;
					out<=5;
				end
			end
			5326: begin
				if(in == 0) begin
					state<=5337;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=1448;
					out<=8;
				end
				if(in == 3) begin
					state<=7269;
					out<=9;
				end
				if(in == 4) begin
					state<=3380;
					out<=10;
				end
			end
			5327: begin
				if(in == 0) begin
					state<=5338;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=1449;
					out<=13;
				end
				if(in == 3) begin
					state<=7270;
					out<=14;
				end
				if(in == 4) begin
					state<=3381;
					out<=15;
				end
			end
			5328: begin
				if(in == 0) begin
					state<=5339;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=1450;
					out<=18;
				end
				if(in == 3) begin
					state<=7271;
					out<=19;
				end
				if(in == 4) begin
					state<=3382;
					out<=20;
				end
			end
			5329: begin
				if(in == 0) begin
					state<=5340;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=1451;
					out<=23;
				end
				if(in == 3) begin
					state<=7272;
					out<=24;
				end
				if(in == 4) begin
					state<=3383;
					out<=25;
				end
			end
			5330: begin
				if(in == 0) begin
					state<=5331;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=1442;
					out<=28;
				end
				if(in == 3) begin
					state<=7263;
					out<=29;
				end
				if(in == 4) begin
					state<=3374;
					out<=30;
				end
			end
			5331: begin
				if(in == 0) begin
					state<=4156;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=258;
					out<=33;
				end
				if(in == 3) begin
					state<=6145;
					out<=34;
				end
				if(in == 4) begin
					state<=2256;
					out<=35;
				end
			end
			5332: begin
				if(in == 0) begin
					state<=4157;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=259;
					out<=38;
				end
				if(in == 3) begin
					state<=6146;
					out<=39;
				end
				if(in == 4) begin
					state<=2257;
					out<=40;
				end
			end
			5333: begin
				if(in == 0) begin
					state<=4158;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=260;
					out<=43;
				end
				if(in == 3) begin
					state<=6147;
					out<=44;
				end
				if(in == 4) begin
					state<=2258;
					out<=45;
				end
			end
			5334: begin
				if(in == 0) begin
					state<=4159;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=261;
					out<=48;
				end
				if(in == 3) begin
					state<=6148;
					out<=49;
				end
				if(in == 4) begin
					state<=2259;
					out<=50;
				end
			end
			5335: begin
				if(in == 0) begin
					state<=4160;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=262;
					out<=53;
				end
				if(in == 3) begin
					state<=6149;
					out<=54;
				end
				if(in == 4) begin
					state<=2260;
					out<=55;
				end
			end
			5336: begin
				if(in == 0) begin
					state<=4161;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=263;
					out<=58;
				end
				if(in == 3) begin
					state<=6150;
					out<=59;
				end
				if(in == 4) begin
					state<=2261;
					out<=60;
				end
			end
			5337: begin
				if(in == 0) begin
					state<=4162;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=264;
					out<=63;
				end
				if(in == 3) begin
					state<=6151;
					out<=64;
				end
				if(in == 4) begin
					state<=2262;
					out<=65;
				end
			end
			5338: begin
				if(in == 0) begin
					state<=4163;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=265;
					out<=68;
				end
				if(in == 3) begin
					state<=6152;
					out<=69;
				end
				if(in == 4) begin
					state<=2263;
					out<=70;
				end
			end
			5339: begin
				if(in == 0) begin
					state<=4164;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=266;
					out<=73;
				end
				if(in == 3) begin
					state<=6153;
					out<=74;
				end
				if(in == 4) begin
					state<=2264;
					out<=75;
				end
			end
			5340: begin
				if(in == 0) begin
					state<=5341;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=1452;
					out<=78;
				end
				if(in == 3) begin
					state<=7273;
					out<=79;
				end
				if(in == 4) begin
					state<=3384;
					out<=80;
				end
			end
			5341: begin
				if(in == 0) begin
					state<=4166;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=268;
					out<=83;
				end
				if(in == 3) begin
					state<=6155;
					out<=84;
				end
				if(in == 4) begin
					state<=2266;
					out<=85;
				end
			end
			5342: begin
				if(in == 0) begin
					state<=5353;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=1464;
					out<=88;
				end
				if(in == 3) begin
					state<=6798;
					out<=89;
				end
				if(in == 4) begin
					state<=2909;
					out<=90;
				end
			end
			5343: begin
				if(in == 0) begin
					state<=5354;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=1465;
					out<=93;
				end
				if(in == 3) begin
					state<=6799;
					out<=94;
				end
				if(in == 4) begin
					state<=2910;
					out<=95;
				end
			end
			5344: begin
				if(in == 0) begin
					state<=5355;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=1466;
					out<=98;
				end
				if(in == 3) begin
					state<=6800;
					out<=99;
				end
				if(in == 4) begin
					state<=2911;
					out<=100;
				end
			end
			5345: begin
				if(in == 0) begin
					state<=5356;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=1467;
					out<=103;
				end
				if(in == 3) begin
					state<=6801;
					out<=104;
				end
				if(in == 4) begin
					state<=2912;
					out<=105;
				end
			end
			5346: begin
				if(in == 0) begin
					state<=5357;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=1468;
					out<=108;
				end
				if(in == 3) begin
					state<=6802;
					out<=109;
				end
				if(in == 4) begin
					state<=2913;
					out<=110;
				end
			end
			5347: begin
				if(in == 0) begin
					state<=5358;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=1469;
					out<=113;
				end
				if(in == 3) begin
					state<=6803;
					out<=114;
				end
				if(in == 4) begin
					state<=2914;
					out<=115;
				end
			end
			5348: begin
				if(in == 0) begin
					state<=5359;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=1470;
					out<=118;
				end
				if(in == 3) begin
					state<=6804;
					out<=119;
				end
				if(in == 4) begin
					state<=2915;
					out<=120;
				end
			end
			5349: begin
				if(in == 0) begin
					state<=5360;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=1471;
					out<=123;
				end
				if(in == 3) begin
					state<=6805;
					out<=124;
				end
				if(in == 4) begin
					state<=2916;
					out<=125;
				end
			end
			5350: begin
				if(in == 0) begin
					state<=5361;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=1472;
					out<=128;
				end
				if(in == 3) begin
					state<=6806;
					out<=129;
				end
				if(in == 4) begin
					state<=2917;
					out<=130;
				end
			end
			5351: begin
				if(in == 0) begin
					state<=5352;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=1463;
					out<=133;
				end
				if(in == 3) begin
					state<=6797;
					out<=134;
				end
				if(in == 4) begin
					state<=2908;
					out<=135;
				end
			end
			5352: begin
				if(in == 0) begin
					state<=5363;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=1474;
					out<=138;
				end
				if(in == 3) begin
					state<=6808;
					out<=139;
				end
				if(in == 4) begin
					state<=2919;
					out<=140;
				end
			end
			5353: begin
				if(in == 0) begin
					state<=5364;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=1475;
					out<=143;
				end
				if(in == 3) begin
					state<=6809;
					out<=144;
				end
				if(in == 4) begin
					state<=2920;
					out<=145;
				end
			end
			5354: begin
				if(in == 0) begin
					state<=5365;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=1476;
					out<=148;
				end
				if(in == 3) begin
					state<=6810;
					out<=149;
				end
				if(in == 4) begin
					state<=2921;
					out<=150;
				end
			end
			5355: begin
				if(in == 0) begin
					state<=5366;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=1477;
					out<=153;
				end
				if(in == 3) begin
					state<=6811;
					out<=154;
				end
				if(in == 4) begin
					state<=2922;
					out<=155;
				end
			end
			5356: begin
				if(in == 0) begin
					state<=5367;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=1478;
					out<=158;
				end
				if(in == 3) begin
					state<=6812;
					out<=159;
				end
				if(in == 4) begin
					state<=2923;
					out<=160;
				end
			end
			5357: begin
				if(in == 0) begin
					state<=5368;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=1479;
					out<=163;
				end
				if(in == 3) begin
					state<=6813;
					out<=164;
				end
				if(in == 4) begin
					state<=2924;
					out<=165;
				end
			end
			5358: begin
				if(in == 0) begin
					state<=5369;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=1480;
					out<=168;
				end
				if(in == 3) begin
					state<=6814;
					out<=169;
				end
				if(in == 4) begin
					state<=2925;
					out<=170;
				end
			end
			5359: begin
				if(in == 0) begin
					state<=5370;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=1481;
					out<=173;
				end
				if(in == 3) begin
					state<=6815;
					out<=174;
				end
				if(in == 4) begin
					state<=2926;
					out<=175;
				end
			end
			5360: begin
				if(in == 0) begin
					state<=5371;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=1482;
					out<=178;
				end
				if(in == 3) begin
					state<=6816;
					out<=179;
				end
				if(in == 4) begin
					state<=2927;
					out<=180;
				end
			end
			5361: begin
				if(in == 0) begin
					state<=5362;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=1473;
					out<=183;
				end
				if(in == 3) begin
					state<=6807;
					out<=184;
				end
				if(in == 4) begin
					state<=2918;
					out<=185;
				end
			end
			5362: begin
				if(in == 0) begin
					state<=4225;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=327;
					out<=188;
				end
				if(in == 3) begin
					state<=6214;
					out<=189;
				end
				if(in == 4) begin
					state<=2325;
					out<=190;
				end
			end
			5363: begin
				if(in == 0) begin
					state<=4226;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=328;
					out<=193;
				end
				if(in == 3) begin
					state<=6215;
					out<=194;
				end
				if(in == 4) begin
					state<=2326;
					out<=195;
				end
			end
			5364: begin
				if(in == 0) begin
					state<=4227;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=329;
					out<=198;
				end
				if(in == 3) begin
					state<=6216;
					out<=199;
				end
				if(in == 4) begin
					state<=2327;
					out<=200;
				end
			end
			5365: begin
				if(in == 0) begin
					state<=4228;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=330;
					out<=203;
				end
				if(in == 3) begin
					state<=6217;
					out<=204;
				end
				if(in == 4) begin
					state<=2328;
					out<=205;
				end
			end
			5366: begin
				if(in == 0) begin
					state<=4229;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=331;
					out<=208;
				end
				if(in == 3) begin
					state<=6218;
					out<=209;
				end
				if(in == 4) begin
					state<=2329;
					out<=210;
				end
			end
			5367: begin
				if(in == 0) begin
					state<=4230;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=332;
					out<=213;
				end
				if(in == 3) begin
					state<=6219;
					out<=214;
				end
				if(in == 4) begin
					state<=2330;
					out<=215;
				end
			end
			5368: begin
				if(in == 0) begin
					state<=4231;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=333;
					out<=218;
				end
				if(in == 3) begin
					state<=6220;
					out<=219;
				end
				if(in == 4) begin
					state<=2331;
					out<=220;
				end
			end
			5369: begin
				if(in == 0) begin
					state<=4232;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=334;
					out<=223;
				end
				if(in == 3) begin
					state<=6221;
					out<=224;
				end
				if(in == 4) begin
					state<=2332;
					out<=225;
				end
			end
			5370: begin
				if(in == 0) begin
					state<=4233;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=335;
					out<=228;
				end
				if(in == 3) begin
					state<=6222;
					out<=229;
				end
				if(in == 4) begin
					state<=2333;
					out<=230;
				end
			end
			5371: begin
				if(in == 0) begin
					state<=5372;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=1483;
					out<=233;
				end
				if(in == 3) begin
					state<=6817;
					out<=234;
				end
				if(in == 4) begin
					state<=2928;
					out<=235;
				end
			end
			5372: begin
				if(in == 0) begin
					state<=4235;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=337;
					out<=238;
				end
				if(in == 3) begin
					state<=6224;
					out<=239;
				end
				if(in == 4) begin
					state<=2335;
					out<=240;
				end
			end
			5373: begin
				if(in == 0) begin
					state<=5384;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=1495;
					out<=243;
				end
				if(in == 3) begin
					state<=7316;
					out<=244;
				end
				if(in == 4) begin
					state<=3427;
					out<=245;
				end
			end
			5374: begin
				if(in == 0) begin
					state<=5385;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=1496;
					out<=248;
				end
				if(in == 3) begin
					state<=7317;
					out<=249;
				end
				if(in == 4) begin
					state<=3428;
					out<=250;
				end
			end
			5375: begin
				if(in == 0) begin
					state<=5386;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=1497;
					out<=253;
				end
				if(in == 3) begin
					state<=7318;
					out<=254;
				end
				if(in == 4) begin
					state<=3429;
					out<=255;
				end
			end
			5376: begin
				if(in == 0) begin
					state<=5387;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=1498;
					out<=2;
				end
				if(in == 3) begin
					state<=7319;
					out<=3;
				end
				if(in == 4) begin
					state<=3430;
					out<=4;
				end
			end
			5377: begin
				if(in == 0) begin
					state<=5388;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=1499;
					out<=7;
				end
				if(in == 3) begin
					state<=7320;
					out<=8;
				end
				if(in == 4) begin
					state<=3431;
					out<=9;
				end
			end
			5378: begin
				if(in == 0) begin
					state<=5389;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=1500;
					out<=12;
				end
				if(in == 3) begin
					state<=7321;
					out<=13;
				end
				if(in == 4) begin
					state<=3432;
					out<=14;
				end
			end
			5379: begin
				if(in == 0) begin
					state<=5390;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=1501;
					out<=17;
				end
				if(in == 3) begin
					state<=7322;
					out<=18;
				end
				if(in == 4) begin
					state<=3433;
					out<=19;
				end
			end
			5380: begin
				if(in == 0) begin
					state<=5391;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=1502;
					out<=22;
				end
				if(in == 3) begin
					state<=7323;
					out<=23;
				end
				if(in == 4) begin
					state<=3434;
					out<=24;
				end
			end
			5381: begin
				if(in == 0) begin
					state<=5392;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=1503;
					out<=27;
				end
				if(in == 3) begin
					state<=7324;
					out<=28;
				end
				if(in == 4) begin
					state<=3435;
					out<=29;
				end
			end
			5382: begin
				if(in == 0) begin
					state<=5383;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=1494;
					out<=32;
				end
				if(in == 3) begin
					state<=7315;
					out<=33;
				end
				if(in == 4) begin
					state<=3426;
					out<=34;
				end
			end
			5383: begin
				if(in == 0) begin
					state<=5394;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=1505;
					out<=37;
				end
				if(in == 3) begin
					state<=7326;
					out<=38;
				end
				if(in == 4) begin
					state<=3437;
					out<=39;
				end
			end
			5384: begin
				if(in == 0) begin
					state<=5395;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=1506;
					out<=42;
				end
				if(in == 3) begin
					state<=7327;
					out<=43;
				end
				if(in == 4) begin
					state<=3438;
					out<=44;
				end
			end
			5385: begin
				if(in == 0) begin
					state<=5396;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=1507;
					out<=47;
				end
				if(in == 3) begin
					state<=7328;
					out<=48;
				end
				if(in == 4) begin
					state<=3439;
					out<=49;
				end
			end
			5386: begin
				if(in == 0) begin
					state<=5397;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=1508;
					out<=52;
				end
				if(in == 3) begin
					state<=7329;
					out<=53;
				end
				if(in == 4) begin
					state<=3440;
					out<=54;
				end
			end
			5387: begin
				if(in == 0) begin
					state<=5398;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=1509;
					out<=57;
				end
				if(in == 3) begin
					state<=7330;
					out<=58;
				end
				if(in == 4) begin
					state<=3441;
					out<=59;
				end
			end
			5388: begin
				if(in == 0) begin
					state<=5399;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=1510;
					out<=62;
				end
				if(in == 3) begin
					state<=7331;
					out<=63;
				end
				if(in == 4) begin
					state<=3442;
					out<=64;
				end
			end
			5389: begin
				if(in == 0) begin
					state<=5400;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=1511;
					out<=67;
				end
				if(in == 3) begin
					state<=7332;
					out<=68;
				end
				if(in == 4) begin
					state<=3443;
					out<=69;
				end
			end
			5390: begin
				if(in == 0) begin
					state<=5401;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=1512;
					out<=72;
				end
				if(in == 3) begin
					state<=7333;
					out<=73;
				end
				if(in == 4) begin
					state<=3444;
					out<=74;
				end
			end
			5391: begin
				if(in == 0) begin
					state<=5402;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=1513;
					out<=77;
				end
				if(in == 3) begin
					state<=7334;
					out<=78;
				end
				if(in == 4) begin
					state<=3445;
					out<=79;
				end
			end
			5392: begin
				if(in == 0) begin
					state<=5393;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=1504;
					out<=82;
				end
				if(in == 3) begin
					state<=7325;
					out<=83;
				end
				if(in == 4) begin
					state<=3436;
					out<=84;
				end
			end
			5393: begin
				if(in == 0) begin
					state<=4363;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=465;
					out<=87;
				end
				if(in == 3) begin
					state<=6352;
					out<=88;
				end
				if(in == 4) begin
					state<=2463;
					out<=89;
				end
			end
			5394: begin
				if(in == 0) begin
					state<=4364;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=466;
					out<=92;
				end
				if(in == 3) begin
					state<=6353;
					out<=93;
				end
				if(in == 4) begin
					state<=2464;
					out<=94;
				end
			end
			5395: begin
				if(in == 0) begin
					state<=4365;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=467;
					out<=97;
				end
				if(in == 3) begin
					state<=6354;
					out<=98;
				end
				if(in == 4) begin
					state<=2465;
					out<=99;
				end
			end
			5396: begin
				if(in == 0) begin
					state<=4366;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=468;
					out<=102;
				end
				if(in == 3) begin
					state<=6355;
					out<=103;
				end
				if(in == 4) begin
					state<=2466;
					out<=104;
				end
			end
			5397: begin
				if(in == 0) begin
					state<=4367;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=469;
					out<=107;
				end
				if(in == 3) begin
					state<=6356;
					out<=108;
				end
				if(in == 4) begin
					state<=2467;
					out<=109;
				end
			end
			5398: begin
				if(in == 0) begin
					state<=4368;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=470;
					out<=112;
				end
				if(in == 3) begin
					state<=6357;
					out<=113;
				end
				if(in == 4) begin
					state<=2468;
					out<=114;
				end
			end
			5399: begin
				if(in == 0) begin
					state<=4369;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=471;
					out<=117;
				end
				if(in == 3) begin
					state<=6358;
					out<=118;
				end
				if(in == 4) begin
					state<=2469;
					out<=119;
				end
			end
			5400: begin
				if(in == 0) begin
					state<=4370;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=472;
					out<=122;
				end
				if(in == 3) begin
					state<=6359;
					out<=123;
				end
				if(in == 4) begin
					state<=2470;
					out<=124;
				end
			end
			5401: begin
				if(in == 0) begin
					state<=4371;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=473;
					out<=127;
				end
				if(in == 3) begin
					state<=6360;
					out<=128;
				end
				if(in == 4) begin
					state<=2471;
					out<=129;
				end
			end
			5402: begin
				if(in == 0) begin
					state<=5403;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=1514;
					out<=132;
				end
				if(in == 3) begin
					state<=7335;
					out<=133;
				end
				if(in == 4) begin
					state<=3446;
					out<=134;
				end
			end
			5403: begin
				if(in == 0) begin
					state<=4373;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=475;
					out<=137;
				end
				if(in == 3) begin
					state<=6362;
					out<=138;
				end
				if(in == 4) begin
					state<=2473;
					out<=139;
				end
			end
			5404: begin
				if(in == 0) begin
					state<=5415;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=1526;
					out<=142;
				end
				if(in == 3) begin
					state<=7347;
					out<=143;
				end
				if(in == 4) begin
					state<=3458;
					out<=144;
				end
			end
			5405: begin
				if(in == 0) begin
					state<=5416;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=1527;
					out<=147;
				end
				if(in == 3) begin
					state<=7348;
					out<=148;
				end
				if(in == 4) begin
					state<=3459;
					out<=149;
				end
			end
			5406: begin
				if(in == 0) begin
					state<=5417;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=1528;
					out<=152;
				end
				if(in == 3) begin
					state<=7349;
					out<=153;
				end
				if(in == 4) begin
					state<=3460;
					out<=154;
				end
			end
			5407: begin
				if(in == 0) begin
					state<=5418;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=1529;
					out<=157;
				end
				if(in == 3) begin
					state<=7350;
					out<=158;
				end
				if(in == 4) begin
					state<=3461;
					out<=159;
				end
			end
			5408: begin
				if(in == 0) begin
					state<=5419;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=1530;
					out<=162;
				end
				if(in == 3) begin
					state<=7351;
					out<=163;
				end
				if(in == 4) begin
					state<=3462;
					out<=164;
				end
			end
			5409: begin
				if(in == 0) begin
					state<=5420;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=1531;
					out<=167;
				end
				if(in == 3) begin
					state<=7352;
					out<=168;
				end
				if(in == 4) begin
					state<=3463;
					out<=169;
				end
			end
			5410: begin
				if(in == 0) begin
					state<=5421;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=1532;
					out<=172;
				end
				if(in == 3) begin
					state<=7353;
					out<=173;
				end
				if(in == 4) begin
					state<=3464;
					out<=174;
				end
			end
			5411: begin
				if(in == 0) begin
					state<=5422;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=1533;
					out<=177;
				end
				if(in == 3) begin
					state<=7354;
					out<=178;
				end
				if(in == 4) begin
					state<=3465;
					out<=179;
				end
			end
			5412: begin
				if(in == 0) begin
					state<=5423;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=1534;
					out<=182;
				end
				if(in == 3) begin
					state<=7355;
					out<=183;
				end
				if(in == 4) begin
					state<=3466;
					out<=184;
				end
			end
			5413: begin
				if(in == 0) begin
					state<=5414;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=1525;
					out<=187;
				end
				if(in == 3) begin
					state<=7346;
					out<=188;
				end
				if(in == 4) begin
					state<=3457;
					out<=189;
				end
			end
			5414: begin
				if(in == 0) begin
					state<=5425;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=1536;
					out<=192;
				end
				if(in == 3) begin
					state<=7357;
					out<=193;
				end
				if(in == 4) begin
					state<=3468;
					out<=194;
				end
			end
			5415: begin
				if(in == 0) begin
					state<=5426;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=1537;
					out<=197;
				end
				if(in == 3) begin
					state<=7358;
					out<=198;
				end
				if(in == 4) begin
					state<=3469;
					out<=199;
				end
			end
			5416: begin
				if(in == 0) begin
					state<=5427;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=1538;
					out<=202;
				end
				if(in == 3) begin
					state<=7359;
					out<=203;
				end
				if(in == 4) begin
					state<=3470;
					out<=204;
				end
			end
			5417: begin
				if(in == 0) begin
					state<=5428;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=1539;
					out<=207;
				end
				if(in == 3) begin
					state<=7360;
					out<=208;
				end
				if(in == 4) begin
					state<=3471;
					out<=209;
				end
			end
			5418: begin
				if(in == 0) begin
					state<=5429;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=1540;
					out<=212;
				end
				if(in == 3) begin
					state<=7361;
					out<=213;
				end
				if(in == 4) begin
					state<=3472;
					out<=214;
				end
			end
			5419: begin
				if(in == 0) begin
					state<=5430;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=1541;
					out<=217;
				end
				if(in == 3) begin
					state<=7362;
					out<=218;
				end
				if(in == 4) begin
					state<=3473;
					out<=219;
				end
			end
			5420: begin
				if(in == 0) begin
					state<=5431;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=1542;
					out<=222;
				end
				if(in == 3) begin
					state<=7363;
					out<=223;
				end
				if(in == 4) begin
					state<=3474;
					out<=224;
				end
			end
			5421: begin
				if(in == 0) begin
					state<=5432;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=1543;
					out<=227;
				end
				if(in == 3) begin
					state<=7364;
					out<=228;
				end
				if(in == 4) begin
					state<=3475;
					out<=229;
				end
			end
			5422: begin
				if(in == 0) begin
					state<=5433;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=1544;
					out<=232;
				end
				if(in == 3) begin
					state<=7365;
					out<=233;
				end
				if(in == 4) begin
					state<=3476;
					out<=234;
				end
			end
			5423: begin
				if(in == 0) begin
					state<=5424;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=1535;
					out<=237;
				end
				if(in == 3) begin
					state<=7356;
					out<=238;
				end
				if(in == 4) begin
					state<=3467;
					out<=239;
				end
			end
			5424: begin
				if(in == 0) begin
					state<=4432;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=534;
					out<=242;
				end
				if(in == 3) begin
					state<=6421;
					out<=243;
				end
				if(in == 4) begin
					state<=2532;
					out<=244;
				end
			end
			5425: begin
				if(in == 0) begin
					state<=4433;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=535;
					out<=247;
				end
				if(in == 3) begin
					state<=6422;
					out<=248;
				end
				if(in == 4) begin
					state<=2533;
					out<=249;
				end
			end
			5426: begin
				if(in == 0) begin
					state<=4434;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=536;
					out<=252;
				end
				if(in == 3) begin
					state<=6423;
					out<=253;
				end
				if(in == 4) begin
					state<=2534;
					out<=254;
				end
			end
			5427: begin
				if(in == 0) begin
					state<=4435;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=537;
					out<=1;
				end
				if(in == 3) begin
					state<=6424;
					out<=2;
				end
				if(in == 4) begin
					state<=2535;
					out<=3;
				end
			end
			5428: begin
				if(in == 0) begin
					state<=4436;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=538;
					out<=6;
				end
				if(in == 3) begin
					state<=6425;
					out<=7;
				end
				if(in == 4) begin
					state<=2536;
					out<=8;
				end
			end
			5429: begin
				if(in == 0) begin
					state<=4437;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=539;
					out<=11;
				end
				if(in == 3) begin
					state<=6426;
					out<=12;
				end
				if(in == 4) begin
					state<=2537;
					out<=13;
				end
			end
			5430: begin
				if(in == 0) begin
					state<=4438;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=540;
					out<=16;
				end
				if(in == 3) begin
					state<=6427;
					out<=17;
				end
				if(in == 4) begin
					state<=2538;
					out<=18;
				end
			end
			5431: begin
				if(in == 0) begin
					state<=4439;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=541;
					out<=21;
				end
				if(in == 3) begin
					state<=6428;
					out<=22;
				end
				if(in == 4) begin
					state<=2539;
					out<=23;
				end
			end
			5432: begin
				if(in == 0) begin
					state<=4440;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=542;
					out<=26;
				end
				if(in == 3) begin
					state<=6429;
					out<=27;
				end
				if(in == 4) begin
					state<=2540;
					out<=28;
				end
			end
			5433: begin
				if(in == 0) begin
					state<=5434;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=1545;
					out<=31;
				end
				if(in == 3) begin
					state<=7366;
					out<=32;
				end
				if(in == 4) begin
					state<=3477;
					out<=33;
				end
			end
			5434: begin
				if(in == 0) begin
					state<=4442;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=544;
					out<=36;
				end
				if(in == 3) begin
					state<=6431;
					out<=37;
				end
				if(in == 4) begin
					state<=2542;
					out<=38;
				end
			end
			5435: begin
				if(in == 0) begin
					state<=5446;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=1557;
					out<=41;
				end
				if(in == 3) begin
					state<=7378;
					out<=42;
				end
				if(in == 4) begin
					state<=3489;
					out<=43;
				end
			end
			5436: begin
				if(in == 0) begin
					state<=5447;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=1558;
					out<=46;
				end
				if(in == 3) begin
					state<=7379;
					out<=47;
				end
				if(in == 4) begin
					state<=3490;
					out<=48;
				end
			end
			5437: begin
				if(in == 0) begin
					state<=5448;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=1559;
					out<=51;
				end
				if(in == 3) begin
					state<=7380;
					out<=52;
				end
				if(in == 4) begin
					state<=3491;
					out<=53;
				end
			end
			5438: begin
				if(in == 0) begin
					state<=5449;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=1560;
					out<=56;
				end
				if(in == 3) begin
					state<=7381;
					out<=57;
				end
				if(in == 4) begin
					state<=3492;
					out<=58;
				end
			end
			5439: begin
				if(in == 0) begin
					state<=5450;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=1561;
					out<=61;
				end
				if(in == 3) begin
					state<=7382;
					out<=62;
				end
				if(in == 4) begin
					state<=3493;
					out<=63;
				end
			end
			5440: begin
				if(in == 0) begin
					state<=5451;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=1562;
					out<=66;
				end
				if(in == 3) begin
					state<=7383;
					out<=67;
				end
				if(in == 4) begin
					state<=3494;
					out<=68;
				end
			end
			5441: begin
				if(in == 0) begin
					state<=5452;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=1563;
					out<=71;
				end
				if(in == 3) begin
					state<=7384;
					out<=72;
				end
				if(in == 4) begin
					state<=3495;
					out<=73;
				end
			end
			5442: begin
				if(in == 0) begin
					state<=5453;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=1564;
					out<=76;
				end
				if(in == 3) begin
					state<=7385;
					out<=77;
				end
				if(in == 4) begin
					state<=3496;
					out<=78;
				end
			end
			5443: begin
				if(in == 0) begin
					state<=5454;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=1565;
					out<=81;
				end
				if(in == 3) begin
					state<=7386;
					out<=82;
				end
				if(in == 4) begin
					state<=3497;
					out<=83;
				end
			end
			5444: begin
				if(in == 0) begin
					state<=5445;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=1556;
					out<=86;
				end
				if(in == 3) begin
					state<=7377;
					out<=87;
				end
				if(in == 4) begin
					state<=3488;
					out<=88;
				end
			end
			5445: begin
				if(in == 0) begin
					state<=5456;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=1567;
					out<=91;
				end
				if(in == 3) begin
					state<=7388;
					out<=92;
				end
				if(in == 4) begin
					state<=3499;
					out<=93;
				end
			end
			5446: begin
				if(in == 0) begin
					state<=5457;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=1568;
					out<=96;
				end
				if(in == 3) begin
					state<=7389;
					out<=97;
				end
				if(in == 4) begin
					state<=3500;
					out<=98;
				end
			end
			5447: begin
				if(in == 0) begin
					state<=5458;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=1569;
					out<=101;
				end
				if(in == 3) begin
					state<=7390;
					out<=102;
				end
				if(in == 4) begin
					state<=3501;
					out<=103;
				end
			end
			5448: begin
				if(in == 0) begin
					state<=5459;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=1570;
					out<=106;
				end
				if(in == 3) begin
					state<=7391;
					out<=107;
				end
				if(in == 4) begin
					state<=3502;
					out<=108;
				end
			end
			5449: begin
				if(in == 0) begin
					state<=5460;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=1571;
					out<=111;
				end
				if(in == 3) begin
					state<=7392;
					out<=112;
				end
				if(in == 4) begin
					state<=3503;
					out<=113;
				end
			end
			5450: begin
				if(in == 0) begin
					state<=5461;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=1572;
					out<=116;
				end
				if(in == 3) begin
					state<=7393;
					out<=117;
				end
				if(in == 4) begin
					state<=3504;
					out<=118;
				end
			end
			5451: begin
				if(in == 0) begin
					state<=5462;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=1573;
					out<=121;
				end
				if(in == 3) begin
					state<=7394;
					out<=122;
				end
				if(in == 4) begin
					state<=3505;
					out<=123;
				end
			end
			5452: begin
				if(in == 0) begin
					state<=5463;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=1574;
					out<=126;
				end
				if(in == 3) begin
					state<=7395;
					out<=127;
				end
				if(in == 4) begin
					state<=3506;
					out<=128;
				end
			end
			5453: begin
				if(in == 0) begin
					state<=5464;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=1575;
					out<=131;
				end
				if(in == 3) begin
					state<=7396;
					out<=132;
				end
				if(in == 4) begin
					state<=3507;
					out<=133;
				end
			end
			5454: begin
				if(in == 0) begin
					state<=5455;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=1566;
					out<=136;
				end
				if(in == 3) begin
					state<=7387;
					out<=137;
				end
				if(in == 4) begin
					state<=3498;
					out<=138;
				end
			end
			5455: begin
				if(in == 0) begin
					state<=4501;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=603;
					out<=141;
				end
				if(in == 3) begin
					state<=6490;
					out<=142;
				end
				if(in == 4) begin
					state<=2601;
					out<=143;
				end
			end
			5456: begin
				if(in == 0) begin
					state<=4502;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=604;
					out<=146;
				end
				if(in == 3) begin
					state<=6491;
					out<=147;
				end
				if(in == 4) begin
					state<=2602;
					out<=148;
				end
			end
			5457: begin
				if(in == 0) begin
					state<=4503;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=605;
					out<=151;
				end
				if(in == 3) begin
					state<=6492;
					out<=152;
				end
				if(in == 4) begin
					state<=2603;
					out<=153;
				end
			end
			5458: begin
				if(in == 0) begin
					state<=4504;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=606;
					out<=156;
				end
				if(in == 3) begin
					state<=6493;
					out<=157;
				end
				if(in == 4) begin
					state<=2604;
					out<=158;
				end
			end
			5459: begin
				if(in == 0) begin
					state<=4505;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=607;
					out<=161;
				end
				if(in == 3) begin
					state<=6494;
					out<=162;
				end
				if(in == 4) begin
					state<=2605;
					out<=163;
				end
			end
			5460: begin
				if(in == 0) begin
					state<=4506;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=608;
					out<=166;
				end
				if(in == 3) begin
					state<=6495;
					out<=167;
				end
				if(in == 4) begin
					state<=2606;
					out<=168;
				end
			end
			5461: begin
				if(in == 0) begin
					state<=4507;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=609;
					out<=171;
				end
				if(in == 3) begin
					state<=6496;
					out<=172;
				end
				if(in == 4) begin
					state<=2607;
					out<=173;
				end
			end
			5462: begin
				if(in == 0) begin
					state<=4508;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=610;
					out<=176;
				end
				if(in == 3) begin
					state<=6497;
					out<=177;
				end
				if(in == 4) begin
					state<=2608;
					out<=178;
				end
			end
			5463: begin
				if(in == 0) begin
					state<=4509;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=611;
					out<=181;
				end
				if(in == 3) begin
					state<=6498;
					out<=182;
				end
				if(in == 4) begin
					state<=2609;
					out<=183;
				end
			end
			5464: begin
				if(in == 0) begin
					state<=5465;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=1576;
					out<=186;
				end
				if(in == 3) begin
					state<=7397;
					out<=187;
				end
				if(in == 4) begin
					state<=3508;
					out<=188;
				end
			end
			5465: begin
				if(in == 0) begin
					state<=4511;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=613;
					out<=191;
				end
				if(in == 3) begin
					state<=6500;
					out<=192;
				end
				if(in == 4) begin
					state<=2611;
					out<=193;
				end
			end
			5466: begin
				if(in == 0) begin
					state<=5477;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=1588;
					out<=196;
				end
				if(in == 3) begin
					state<=7130;
					out<=197;
				end
				if(in == 4) begin
					state<=3241;
					out<=198;
				end
			end
			5467: begin
				if(in == 0) begin
					state<=5478;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=1589;
					out<=201;
				end
				if(in == 3) begin
					state<=7131;
					out<=202;
				end
				if(in == 4) begin
					state<=3242;
					out<=203;
				end
			end
			5468: begin
				if(in == 0) begin
					state<=5479;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=1590;
					out<=206;
				end
				if(in == 3) begin
					state<=7132;
					out<=207;
				end
				if(in == 4) begin
					state<=3243;
					out<=208;
				end
			end
			5469: begin
				if(in == 0) begin
					state<=5480;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=1591;
					out<=211;
				end
				if(in == 3) begin
					state<=7133;
					out<=212;
				end
				if(in == 4) begin
					state<=3244;
					out<=213;
				end
			end
			5470: begin
				if(in == 0) begin
					state<=5481;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=1592;
					out<=216;
				end
				if(in == 3) begin
					state<=7134;
					out<=217;
				end
				if(in == 4) begin
					state<=3245;
					out<=218;
				end
			end
			5471: begin
				if(in == 0) begin
					state<=5482;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=1593;
					out<=221;
				end
				if(in == 3) begin
					state<=7135;
					out<=222;
				end
				if(in == 4) begin
					state<=3246;
					out<=223;
				end
			end
			5472: begin
				if(in == 0) begin
					state<=5483;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=1594;
					out<=226;
				end
				if(in == 3) begin
					state<=7136;
					out<=227;
				end
				if(in == 4) begin
					state<=3247;
					out<=228;
				end
			end
			5473: begin
				if(in == 0) begin
					state<=5484;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=1595;
					out<=231;
				end
				if(in == 3) begin
					state<=7137;
					out<=232;
				end
				if(in == 4) begin
					state<=3248;
					out<=233;
				end
			end
			5474: begin
				if(in == 0) begin
					state<=5485;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=1596;
					out<=236;
				end
				if(in == 3) begin
					state<=7138;
					out<=237;
				end
				if(in == 4) begin
					state<=3249;
					out<=238;
				end
			end
			5475: begin
				if(in == 0) begin
					state<=5476;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=1587;
					out<=241;
				end
				if(in == 3) begin
					state<=7129;
					out<=242;
				end
				if(in == 4) begin
					state<=3240;
					out<=243;
				end
			end
			5476: begin
				if(in == 0) begin
					state<=5487;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=1598;
					out<=246;
				end
				if(in == 3) begin
					state<=7140;
					out<=247;
				end
				if(in == 4) begin
					state<=3251;
					out<=248;
				end
			end
			5477: begin
				if(in == 0) begin
					state<=5488;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=1599;
					out<=251;
				end
				if(in == 3) begin
					state<=7141;
					out<=252;
				end
				if(in == 4) begin
					state<=3252;
					out<=253;
				end
			end
			5478: begin
				if(in == 0) begin
					state<=5489;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=1600;
					out<=0;
				end
				if(in == 3) begin
					state<=7142;
					out<=1;
				end
				if(in == 4) begin
					state<=3253;
					out<=2;
				end
			end
			5479: begin
				if(in == 0) begin
					state<=5490;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=1601;
					out<=5;
				end
				if(in == 3) begin
					state<=7143;
					out<=6;
				end
				if(in == 4) begin
					state<=3254;
					out<=7;
				end
			end
			5480: begin
				if(in == 0) begin
					state<=5491;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=1602;
					out<=10;
				end
				if(in == 3) begin
					state<=7144;
					out<=11;
				end
				if(in == 4) begin
					state<=3255;
					out<=12;
				end
			end
			5481: begin
				if(in == 0) begin
					state<=5492;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=1603;
					out<=15;
				end
				if(in == 3) begin
					state<=7145;
					out<=16;
				end
				if(in == 4) begin
					state<=3256;
					out<=17;
				end
			end
			5482: begin
				if(in == 0) begin
					state<=5493;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=1604;
					out<=20;
				end
				if(in == 3) begin
					state<=7146;
					out<=21;
				end
				if(in == 4) begin
					state<=3257;
					out<=22;
				end
			end
			5483: begin
				if(in == 0) begin
					state<=5494;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=1605;
					out<=25;
				end
				if(in == 3) begin
					state<=7147;
					out<=26;
				end
				if(in == 4) begin
					state<=3258;
					out<=27;
				end
			end
			5484: begin
				if(in == 0) begin
					state<=5495;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=1606;
					out<=30;
				end
				if(in == 3) begin
					state<=7148;
					out<=31;
				end
				if(in == 4) begin
					state<=3259;
					out<=32;
				end
			end
			5485: begin
				if(in == 0) begin
					state<=5486;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=1597;
					out<=35;
				end
				if(in == 3) begin
					state<=7139;
					out<=36;
				end
				if(in == 4) begin
					state<=3250;
					out<=37;
				end
			end
			5486: begin
				if(in == 0) begin
					state<=4570;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=672;
					out<=40;
				end
				if(in == 3) begin
					state<=6559;
					out<=41;
				end
				if(in == 4) begin
					state<=2670;
					out<=42;
				end
			end
			5487: begin
				if(in == 0) begin
					state<=4571;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=673;
					out<=45;
				end
				if(in == 3) begin
					state<=6560;
					out<=46;
				end
				if(in == 4) begin
					state<=2671;
					out<=47;
				end
			end
			5488: begin
				if(in == 0) begin
					state<=4572;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=674;
					out<=50;
				end
				if(in == 3) begin
					state<=6561;
					out<=51;
				end
				if(in == 4) begin
					state<=2672;
					out<=52;
				end
			end
			5489: begin
				if(in == 0) begin
					state<=4573;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=675;
					out<=55;
				end
				if(in == 3) begin
					state<=6562;
					out<=56;
				end
				if(in == 4) begin
					state<=2673;
					out<=57;
				end
			end
			5490: begin
				if(in == 0) begin
					state<=4574;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=676;
					out<=60;
				end
				if(in == 3) begin
					state<=6563;
					out<=61;
				end
				if(in == 4) begin
					state<=2674;
					out<=62;
				end
			end
			5491: begin
				if(in == 0) begin
					state<=4575;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=677;
					out<=65;
				end
				if(in == 3) begin
					state<=6564;
					out<=66;
				end
				if(in == 4) begin
					state<=2675;
					out<=67;
				end
			end
			5492: begin
				if(in == 0) begin
					state<=4576;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=678;
					out<=70;
				end
				if(in == 3) begin
					state<=6565;
					out<=71;
				end
				if(in == 4) begin
					state<=2676;
					out<=72;
				end
			end
			5493: begin
				if(in == 0) begin
					state<=4577;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=679;
					out<=75;
				end
				if(in == 3) begin
					state<=6566;
					out<=76;
				end
				if(in == 4) begin
					state<=2677;
					out<=77;
				end
			end
			5494: begin
				if(in == 0) begin
					state<=4578;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=680;
					out<=80;
				end
				if(in == 3) begin
					state<=6567;
					out<=81;
				end
				if(in == 4) begin
					state<=2678;
					out<=82;
				end
			end
			5495: begin
				if(in == 0) begin
					state<=5496;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=1607;
					out<=85;
				end
				if(in == 3) begin
					state<=7149;
					out<=86;
				end
				if(in == 4) begin
					state<=3260;
					out<=87;
				end
			end
			5496: begin
				if(in == 0) begin
					state<=4580;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=682;
					out<=90;
				end
				if(in == 3) begin
					state<=6569;
					out<=91;
				end
				if(in == 4) begin
					state<=2680;
					out<=92;
				end
			end
			5497: begin
				if(in == 0) begin
					state<=5508;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=1619;
					out<=95;
				end
				if(in == 3) begin
					state<=7409;
					out<=96;
				end
				if(in == 4) begin
					state<=3520;
					out<=97;
				end
			end
			5498: begin
				if(in == 0) begin
					state<=5509;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=1620;
					out<=100;
				end
				if(in == 3) begin
					state<=7410;
					out<=101;
				end
				if(in == 4) begin
					state<=3521;
					out<=102;
				end
			end
			5499: begin
				if(in == 0) begin
					state<=5510;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=1621;
					out<=105;
				end
				if(in == 3) begin
					state<=7411;
					out<=106;
				end
				if(in == 4) begin
					state<=3522;
					out<=107;
				end
			end
			5500: begin
				if(in == 0) begin
					state<=5511;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=1622;
					out<=110;
				end
				if(in == 3) begin
					state<=7412;
					out<=111;
				end
				if(in == 4) begin
					state<=3523;
					out<=112;
				end
			end
			5501: begin
				if(in == 0) begin
					state<=5512;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=1623;
					out<=115;
				end
				if(in == 3) begin
					state<=7413;
					out<=116;
				end
				if(in == 4) begin
					state<=3524;
					out<=117;
				end
			end
			5502: begin
				if(in == 0) begin
					state<=5513;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=1624;
					out<=120;
				end
				if(in == 3) begin
					state<=7414;
					out<=121;
				end
				if(in == 4) begin
					state<=3525;
					out<=122;
				end
			end
			5503: begin
				if(in == 0) begin
					state<=5514;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=1625;
					out<=125;
				end
				if(in == 3) begin
					state<=7415;
					out<=126;
				end
				if(in == 4) begin
					state<=3526;
					out<=127;
				end
			end
			5504: begin
				if(in == 0) begin
					state<=5515;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=1626;
					out<=130;
				end
				if(in == 3) begin
					state<=7416;
					out<=131;
				end
				if(in == 4) begin
					state<=3527;
					out<=132;
				end
			end
			5505: begin
				if(in == 0) begin
					state<=5516;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=1627;
					out<=135;
				end
				if(in == 3) begin
					state<=7417;
					out<=136;
				end
				if(in == 4) begin
					state<=3528;
					out<=137;
				end
			end
			5506: begin
				if(in == 0) begin
					state<=5507;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=1618;
					out<=140;
				end
				if(in == 3) begin
					state<=7408;
					out<=141;
				end
				if(in == 4) begin
					state<=3519;
					out<=142;
				end
			end
			5507: begin
				if(in == 0) begin
					state<=5518;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=1629;
					out<=145;
				end
				if(in == 3) begin
					state<=7419;
					out<=146;
				end
				if(in == 4) begin
					state<=3530;
					out<=147;
				end
			end
			5508: begin
				if(in == 0) begin
					state<=5519;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=1630;
					out<=150;
				end
				if(in == 3) begin
					state<=7420;
					out<=151;
				end
				if(in == 4) begin
					state<=3531;
					out<=152;
				end
			end
			5509: begin
				if(in == 0) begin
					state<=5520;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=1631;
					out<=155;
				end
				if(in == 3) begin
					state<=7421;
					out<=156;
				end
				if(in == 4) begin
					state<=3532;
					out<=157;
				end
			end
			5510: begin
				if(in == 0) begin
					state<=5521;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=1632;
					out<=160;
				end
				if(in == 3) begin
					state<=7422;
					out<=161;
				end
				if(in == 4) begin
					state<=3533;
					out<=162;
				end
			end
			5511: begin
				if(in == 0) begin
					state<=5522;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=1633;
					out<=165;
				end
				if(in == 3) begin
					state<=7423;
					out<=166;
				end
				if(in == 4) begin
					state<=3534;
					out<=167;
				end
			end
			5512: begin
				if(in == 0) begin
					state<=5523;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=1634;
					out<=170;
				end
				if(in == 3) begin
					state<=7424;
					out<=171;
				end
				if(in == 4) begin
					state<=3535;
					out<=172;
				end
			end
			5513: begin
				if(in == 0) begin
					state<=5524;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=1635;
					out<=175;
				end
				if(in == 3) begin
					state<=7425;
					out<=176;
				end
				if(in == 4) begin
					state<=3536;
					out<=177;
				end
			end
			5514: begin
				if(in == 0) begin
					state<=5525;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=1636;
					out<=180;
				end
				if(in == 3) begin
					state<=7426;
					out<=181;
				end
				if(in == 4) begin
					state<=3537;
					out<=182;
				end
			end
			5515: begin
				if(in == 0) begin
					state<=5526;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=1637;
					out<=185;
				end
				if(in == 3) begin
					state<=7427;
					out<=186;
				end
				if(in == 4) begin
					state<=3538;
					out<=187;
				end
			end
			5516: begin
				if(in == 0) begin
					state<=5517;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=1628;
					out<=190;
				end
				if(in == 3) begin
					state<=7418;
					out<=191;
				end
				if(in == 4) begin
					state<=3529;
					out<=192;
				end
			end
			5517: begin
				if(in == 0) begin
					state<=5528;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=1639;
					out<=195;
				end
				if(in == 3) begin
					state<=7429;
					out<=196;
				end
				if(in == 4) begin
					state<=3540;
					out<=197;
				end
			end
			5518: begin
				if(in == 0) begin
					state<=5529;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=1640;
					out<=200;
				end
				if(in == 3) begin
					state<=7430;
					out<=201;
				end
				if(in == 4) begin
					state<=3541;
					out<=202;
				end
			end
			5519: begin
				if(in == 0) begin
					state<=5530;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=1641;
					out<=205;
				end
				if(in == 3) begin
					state<=7431;
					out<=206;
				end
				if(in == 4) begin
					state<=3542;
					out<=207;
				end
			end
			5520: begin
				if(in == 0) begin
					state<=5531;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=1642;
					out<=210;
				end
				if(in == 3) begin
					state<=7432;
					out<=211;
				end
				if(in == 4) begin
					state<=3543;
					out<=212;
				end
			end
			5521: begin
				if(in == 0) begin
					state<=5532;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=1643;
					out<=215;
				end
				if(in == 3) begin
					state<=7433;
					out<=216;
				end
				if(in == 4) begin
					state<=3544;
					out<=217;
				end
			end
			5522: begin
				if(in == 0) begin
					state<=5533;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=1644;
					out<=220;
				end
				if(in == 3) begin
					state<=7434;
					out<=221;
				end
				if(in == 4) begin
					state<=3545;
					out<=222;
				end
			end
			5523: begin
				if(in == 0) begin
					state<=5534;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=1645;
					out<=225;
				end
				if(in == 3) begin
					state<=7435;
					out<=226;
				end
				if(in == 4) begin
					state<=3546;
					out<=227;
				end
			end
			5524: begin
				if(in == 0) begin
					state<=5535;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=1646;
					out<=230;
				end
				if(in == 3) begin
					state<=7436;
					out<=231;
				end
				if(in == 4) begin
					state<=3547;
					out<=232;
				end
			end
			5525: begin
				if(in == 0) begin
					state<=5536;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=1647;
					out<=235;
				end
				if(in == 3) begin
					state<=7437;
					out<=236;
				end
				if(in == 4) begin
					state<=3548;
					out<=237;
				end
			end
			5526: begin
				if(in == 0) begin
					state<=5527;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=1638;
					out<=240;
				end
				if(in == 3) begin
					state<=7428;
					out<=241;
				end
				if(in == 4) begin
					state<=3539;
					out<=242;
				end
			end
			5527: begin
				if(in == 0) begin
					state<=5538;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=1649;
					out<=245;
				end
				if(in == 3) begin
					state<=7439;
					out<=246;
				end
				if(in == 4) begin
					state<=3550;
					out<=247;
				end
			end
			5528: begin
				if(in == 0) begin
					state<=5539;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=1650;
					out<=250;
				end
				if(in == 3) begin
					state<=7440;
					out<=251;
				end
				if(in == 4) begin
					state<=3551;
					out<=252;
				end
			end
			5529: begin
				if(in == 0) begin
					state<=5540;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=1651;
					out<=255;
				end
				if(in == 3) begin
					state<=7441;
					out<=0;
				end
				if(in == 4) begin
					state<=3552;
					out<=1;
				end
			end
			5530: begin
				if(in == 0) begin
					state<=5541;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=1652;
					out<=4;
				end
				if(in == 3) begin
					state<=7442;
					out<=5;
				end
				if(in == 4) begin
					state<=3553;
					out<=6;
				end
			end
			5531: begin
				if(in == 0) begin
					state<=5542;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=1653;
					out<=9;
				end
				if(in == 3) begin
					state<=7443;
					out<=10;
				end
				if(in == 4) begin
					state<=3554;
					out<=11;
				end
			end
			5532: begin
				if(in == 0) begin
					state<=5543;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=1654;
					out<=14;
				end
				if(in == 3) begin
					state<=7444;
					out<=15;
				end
				if(in == 4) begin
					state<=3555;
					out<=16;
				end
			end
			5533: begin
				if(in == 0) begin
					state<=5544;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=1655;
					out<=19;
				end
				if(in == 3) begin
					state<=7445;
					out<=20;
				end
				if(in == 4) begin
					state<=3556;
					out<=21;
				end
			end
			5534: begin
				if(in == 0) begin
					state<=5545;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=1656;
					out<=24;
				end
				if(in == 3) begin
					state<=7446;
					out<=25;
				end
				if(in == 4) begin
					state<=3557;
					out<=26;
				end
			end
			5535: begin
				if(in == 0) begin
					state<=5546;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=1657;
					out<=29;
				end
				if(in == 3) begin
					state<=7447;
					out<=30;
				end
				if(in == 4) begin
					state<=3558;
					out<=31;
				end
			end
			5536: begin
				if(in == 0) begin
					state<=5537;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=1648;
					out<=34;
				end
				if(in == 3) begin
					state<=7438;
					out<=35;
				end
				if(in == 4) begin
					state<=3549;
					out<=36;
				end
			end
			5537: begin
				if(in == 0) begin
					state<=5548;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=1659;
					out<=39;
				end
				if(in == 3) begin
					state<=7449;
					out<=40;
				end
				if(in == 4) begin
					state<=3560;
					out<=41;
				end
			end
			5538: begin
				if(in == 0) begin
					state<=5549;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=1660;
					out<=44;
				end
				if(in == 3) begin
					state<=7450;
					out<=45;
				end
				if(in == 4) begin
					state<=3561;
					out<=46;
				end
			end
			5539: begin
				if(in == 0) begin
					state<=5550;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=1661;
					out<=49;
				end
				if(in == 3) begin
					state<=7451;
					out<=50;
				end
				if(in == 4) begin
					state<=3562;
					out<=51;
				end
			end
			5540: begin
				if(in == 0) begin
					state<=5551;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=1662;
					out<=54;
				end
				if(in == 3) begin
					state<=7452;
					out<=55;
				end
				if(in == 4) begin
					state<=3563;
					out<=56;
				end
			end
			5541: begin
				if(in == 0) begin
					state<=5552;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=1663;
					out<=59;
				end
				if(in == 3) begin
					state<=7453;
					out<=60;
				end
				if(in == 4) begin
					state<=3564;
					out<=61;
				end
			end
			5542: begin
				if(in == 0) begin
					state<=5553;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=1664;
					out<=64;
				end
				if(in == 3) begin
					state<=7454;
					out<=65;
				end
				if(in == 4) begin
					state<=3565;
					out<=66;
				end
			end
			5543: begin
				if(in == 0) begin
					state<=5554;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=1665;
					out<=69;
				end
				if(in == 3) begin
					state<=7455;
					out<=70;
				end
				if(in == 4) begin
					state<=3566;
					out<=71;
				end
			end
			5544: begin
				if(in == 0) begin
					state<=5555;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=1666;
					out<=74;
				end
				if(in == 3) begin
					state<=7456;
					out<=75;
				end
				if(in == 4) begin
					state<=3567;
					out<=76;
				end
			end
			5545: begin
				if(in == 0) begin
					state<=5556;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=1667;
					out<=79;
				end
				if(in == 3) begin
					state<=7457;
					out<=80;
				end
				if(in == 4) begin
					state<=3568;
					out<=81;
				end
			end
			5546: begin
				if(in == 0) begin
					state<=5547;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=1658;
					out<=84;
				end
				if(in == 3) begin
					state<=7448;
					out<=85;
				end
				if(in == 4) begin
					state<=3559;
					out<=86;
				end
			end
			5547: begin
				if(in == 0) begin
					state<=5558;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=1669;
					out<=89;
				end
				if(in == 3) begin
					state<=7459;
					out<=90;
				end
				if(in == 4) begin
					state<=3570;
					out<=91;
				end
			end
			5548: begin
				if(in == 0) begin
					state<=5559;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=1670;
					out<=94;
				end
				if(in == 3) begin
					state<=7460;
					out<=95;
				end
				if(in == 4) begin
					state<=3571;
					out<=96;
				end
			end
			5549: begin
				if(in == 0) begin
					state<=5560;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=1671;
					out<=99;
				end
				if(in == 3) begin
					state<=7461;
					out<=100;
				end
				if(in == 4) begin
					state<=3572;
					out<=101;
				end
			end
			5550: begin
				if(in == 0) begin
					state<=5561;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=1672;
					out<=104;
				end
				if(in == 3) begin
					state<=7462;
					out<=105;
				end
				if(in == 4) begin
					state<=3573;
					out<=106;
				end
			end
			5551: begin
				if(in == 0) begin
					state<=5562;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=1673;
					out<=109;
				end
				if(in == 3) begin
					state<=7463;
					out<=110;
				end
				if(in == 4) begin
					state<=3574;
					out<=111;
				end
			end
			5552: begin
				if(in == 0) begin
					state<=5563;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=1674;
					out<=114;
				end
				if(in == 3) begin
					state<=7464;
					out<=115;
				end
				if(in == 4) begin
					state<=3575;
					out<=116;
				end
			end
			5553: begin
				if(in == 0) begin
					state<=5564;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=1675;
					out<=119;
				end
				if(in == 3) begin
					state<=7465;
					out<=120;
				end
				if(in == 4) begin
					state<=3576;
					out<=121;
				end
			end
			5554: begin
				if(in == 0) begin
					state<=5565;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=1676;
					out<=124;
				end
				if(in == 3) begin
					state<=7466;
					out<=125;
				end
				if(in == 4) begin
					state<=3577;
					out<=126;
				end
			end
			5555: begin
				if(in == 0) begin
					state<=5566;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=1677;
					out<=129;
				end
				if(in == 3) begin
					state<=7467;
					out<=130;
				end
				if(in == 4) begin
					state<=3578;
					out<=131;
				end
			end
			5556: begin
				if(in == 0) begin
					state<=5557;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=1668;
					out<=134;
				end
				if(in == 3) begin
					state<=7458;
					out<=135;
				end
				if(in == 4) begin
					state<=3569;
					out<=136;
				end
			end
			5557: begin
				if(in == 0) begin
					state<=5568;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=1679;
					out<=139;
				end
				if(in == 3) begin
					state<=7469;
					out<=140;
				end
				if(in == 4) begin
					state<=3580;
					out<=141;
				end
			end
			5558: begin
				if(in == 0) begin
					state<=5569;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=1680;
					out<=144;
				end
				if(in == 3) begin
					state<=7470;
					out<=145;
				end
				if(in == 4) begin
					state<=3581;
					out<=146;
				end
			end
			5559: begin
				if(in == 0) begin
					state<=5570;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=1681;
					out<=149;
				end
				if(in == 3) begin
					state<=7471;
					out<=150;
				end
				if(in == 4) begin
					state<=3582;
					out<=151;
				end
			end
			5560: begin
				if(in == 0) begin
					state<=5571;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=1682;
					out<=154;
				end
				if(in == 3) begin
					state<=7472;
					out<=155;
				end
				if(in == 4) begin
					state<=3583;
					out<=156;
				end
			end
			5561: begin
				if(in == 0) begin
					state<=5572;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=1683;
					out<=159;
				end
				if(in == 3) begin
					state<=7473;
					out<=160;
				end
				if(in == 4) begin
					state<=3584;
					out<=161;
				end
			end
			5562: begin
				if(in == 0) begin
					state<=5573;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=1684;
					out<=164;
				end
				if(in == 3) begin
					state<=7474;
					out<=165;
				end
				if(in == 4) begin
					state<=3585;
					out<=166;
				end
			end
			5563: begin
				if(in == 0) begin
					state<=5574;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=1685;
					out<=169;
				end
				if(in == 3) begin
					state<=7475;
					out<=170;
				end
				if(in == 4) begin
					state<=3586;
					out<=171;
				end
			end
			5564: begin
				if(in == 0) begin
					state<=5575;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=1686;
					out<=174;
				end
				if(in == 3) begin
					state<=7476;
					out<=175;
				end
				if(in == 4) begin
					state<=3587;
					out<=176;
				end
			end
			5565: begin
				if(in == 0) begin
					state<=5576;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=1687;
					out<=179;
				end
				if(in == 3) begin
					state<=7477;
					out<=180;
				end
				if(in == 4) begin
					state<=3588;
					out<=181;
				end
			end
			5566: begin
				if(in == 0) begin
					state<=5567;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=1678;
					out<=184;
				end
				if(in == 3) begin
					state<=7468;
					out<=185;
				end
				if(in == 4) begin
					state<=3579;
					out<=186;
				end
			end
			5567: begin
				if(in == 0) begin
					state<=5578;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=1689;
					out<=189;
				end
				if(in == 3) begin
					state<=7479;
					out<=190;
				end
				if(in == 4) begin
					state<=3590;
					out<=191;
				end
			end
			5568: begin
				if(in == 0) begin
					state<=5579;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=1690;
					out<=194;
				end
				if(in == 3) begin
					state<=7480;
					out<=195;
				end
				if(in == 4) begin
					state<=3591;
					out<=196;
				end
			end
			5569: begin
				if(in == 0) begin
					state<=5580;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=1691;
					out<=199;
				end
				if(in == 3) begin
					state<=7481;
					out<=200;
				end
				if(in == 4) begin
					state<=3592;
					out<=201;
				end
			end
			5570: begin
				if(in == 0) begin
					state<=5581;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=1692;
					out<=204;
				end
				if(in == 3) begin
					state<=7482;
					out<=205;
				end
				if(in == 4) begin
					state<=3593;
					out<=206;
				end
			end
			5571: begin
				if(in == 0) begin
					state<=5582;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=1693;
					out<=209;
				end
				if(in == 3) begin
					state<=7483;
					out<=210;
				end
				if(in == 4) begin
					state<=3594;
					out<=211;
				end
			end
			5572: begin
				if(in == 0) begin
					state<=5583;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=1694;
					out<=214;
				end
				if(in == 3) begin
					state<=7484;
					out<=215;
				end
				if(in == 4) begin
					state<=3595;
					out<=216;
				end
			end
			5573: begin
				if(in == 0) begin
					state<=5584;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=1695;
					out<=219;
				end
				if(in == 3) begin
					state<=7485;
					out<=220;
				end
				if(in == 4) begin
					state<=3596;
					out<=221;
				end
			end
			5574: begin
				if(in == 0) begin
					state<=5585;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=1696;
					out<=224;
				end
				if(in == 3) begin
					state<=7486;
					out<=225;
				end
				if(in == 4) begin
					state<=3597;
					out<=226;
				end
			end
			5575: begin
				if(in == 0) begin
					state<=5586;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=1697;
					out<=229;
				end
				if(in == 3) begin
					state<=7487;
					out<=230;
				end
				if(in == 4) begin
					state<=3598;
					out<=231;
				end
			end
			5576: begin
				if(in == 0) begin
					state<=5577;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=1688;
					out<=234;
				end
				if(in == 3) begin
					state<=7478;
					out<=235;
				end
				if(in == 4) begin
					state<=3589;
					out<=236;
				end
			end
			5577: begin
				if(in == 0) begin
					state<=5588;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=1699;
					out<=239;
				end
				if(in == 3) begin
					state<=7489;
					out<=240;
				end
				if(in == 4) begin
					state<=3600;
					out<=241;
				end
			end
			5578: begin
				if(in == 0) begin
					state<=5589;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=1700;
					out<=244;
				end
				if(in == 3) begin
					state<=7490;
					out<=245;
				end
				if(in == 4) begin
					state<=3601;
					out<=246;
				end
			end
			5579: begin
				if(in == 0) begin
					state<=5590;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=1701;
					out<=249;
				end
				if(in == 3) begin
					state<=7491;
					out<=250;
				end
				if(in == 4) begin
					state<=3602;
					out<=251;
				end
			end
			5580: begin
				if(in == 0) begin
					state<=5591;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=1702;
					out<=254;
				end
				if(in == 3) begin
					state<=7492;
					out<=255;
				end
				if(in == 4) begin
					state<=3603;
					out<=0;
				end
			end
			5581: begin
				if(in == 0) begin
					state<=5592;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=1703;
					out<=3;
				end
				if(in == 3) begin
					state<=7493;
					out<=4;
				end
				if(in == 4) begin
					state<=3604;
					out<=5;
				end
			end
			5582: begin
				if(in == 0) begin
					state<=5593;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=1704;
					out<=8;
				end
				if(in == 3) begin
					state<=7494;
					out<=9;
				end
				if(in == 4) begin
					state<=3605;
					out<=10;
				end
			end
			5583: begin
				if(in == 0) begin
					state<=5594;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=1705;
					out<=13;
				end
				if(in == 3) begin
					state<=7495;
					out<=14;
				end
				if(in == 4) begin
					state<=3606;
					out<=15;
				end
			end
			5584: begin
				if(in == 0) begin
					state<=5595;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=1706;
					out<=18;
				end
				if(in == 3) begin
					state<=7496;
					out<=19;
				end
				if(in == 4) begin
					state<=3607;
					out<=20;
				end
			end
			5585: begin
				if(in == 0) begin
					state<=5596;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=1707;
					out<=23;
				end
				if(in == 3) begin
					state<=7497;
					out<=24;
				end
				if(in == 4) begin
					state<=3608;
					out<=25;
				end
			end
			5586: begin
				if(in == 0) begin
					state<=5587;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=1698;
					out<=28;
				end
				if(in == 3) begin
					state<=7488;
					out<=29;
				end
				if(in == 4) begin
					state<=3599;
					out<=30;
				end
			end
			5587: begin
				if(in == 0) begin
					state<=5598;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=1709;
					out<=33;
				end
				if(in == 3) begin
					state<=7499;
					out<=34;
				end
				if(in == 4) begin
					state<=3610;
					out<=35;
				end
			end
			5588: begin
				if(in == 0) begin
					state<=5599;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=1710;
					out<=38;
				end
				if(in == 3) begin
					state<=7500;
					out<=39;
				end
				if(in == 4) begin
					state<=3611;
					out<=40;
				end
			end
			5589: begin
				if(in == 0) begin
					state<=5600;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=1711;
					out<=43;
				end
				if(in == 3) begin
					state<=7501;
					out<=44;
				end
				if(in == 4) begin
					state<=3612;
					out<=45;
				end
			end
			5590: begin
				if(in == 0) begin
					state<=5601;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=1712;
					out<=48;
				end
				if(in == 3) begin
					state<=7502;
					out<=49;
				end
				if(in == 4) begin
					state<=3613;
					out<=50;
				end
			end
			5591: begin
				if(in == 0) begin
					state<=5602;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=1713;
					out<=53;
				end
				if(in == 3) begin
					state<=7503;
					out<=54;
				end
				if(in == 4) begin
					state<=3614;
					out<=55;
				end
			end
			5592: begin
				if(in == 0) begin
					state<=5603;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=1714;
					out<=58;
				end
				if(in == 3) begin
					state<=7504;
					out<=59;
				end
				if(in == 4) begin
					state<=3615;
					out<=60;
				end
			end
			5593: begin
				if(in == 0) begin
					state<=5604;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=1715;
					out<=63;
				end
				if(in == 3) begin
					state<=7505;
					out<=64;
				end
				if(in == 4) begin
					state<=3616;
					out<=65;
				end
			end
			5594: begin
				if(in == 0) begin
					state<=5605;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=1716;
					out<=68;
				end
				if(in == 3) begin
					state<=7506;
					out<=69;
				end
				if(in == 4) begin
					state<=3617;
					out<=70;
				end
			end
			5595: begin
				if(in == 0) begin
					state<=5606;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=1717;
					out<=73;
				end
				if(in == 3) begin
					state<=7507;
					out<=74;
				end
				if(in == 4) begin
					state<=3618;
					out<=75;
				end
			end
			5596: begin
				if(in == 0) begin
					state<=5597;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=1708;
					out<=78;
				end
				if(in == 3) begin
					state<=7498;
					out<=79;
				end
				if(in == 4) begin
					state<=3609;
					out<=80;
				end
			end
			5597: begin
				if(in == 0) begin
					state<=5608;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=1719;
					out<=83;
				end
				if(in == 3) begin
					state<=7509;
					out<=84;
				end
				if(in == 4) begin
					state<=3620;
					out<=85;
				end
			end
			5598: begin
				if(in == 0) begin
					state<=5609;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=1720;
					out<=88;
				end
				if(in == 3) begin
					state<=7510;
					out<=89;
				end
				if(in == 4) begin
					state<=3621;
					out<=90;
				end
			end
			5599: begin
				if(in == 0) begin
					state<=5610;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=1721;
					out<=93;
				end
				if(in == 3) begin
					state<=7511;
					out<=94;
				end
				if(in == 4) begin
					state<=3622;
					out<=95;
				end
			end
			5600: begin
				if(in == 0) begin
					state<=5611;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=1722;
					out<=98;
				end
				if(in == 3) begin
					state<=7512;
					out<=99;
				end
				if(in == 4) begin
					state<=3623;
					out<=100;
				end
			end
			5601: begin
				if(in == 0) begin
					state<=5612;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=1723;
					out<=103;
				end
				if(in == 3) begin
					state<=7513;
					out<=104;
				end
				if(in == 4) begin
					state<=3624;
					out<=105;
				end
			end
			5602: begin
				if(in == 0) begin
					state<=5613;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=1724;
					out<=108;
				end
				if(in == 3) begin
					state<=7514;
					out<=109;
				end
				if(in == 4) begin
					state<=3625;
					out<=110;
				end
			end
			5603: begin
				if(in == 0) begin
					state<=5614;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=1725;
					out<=113;
				end
				if(in == 3) begin
					state<=7515;
					out<=114;
				end
				if(in == 4) begin
					state<=3626;
					out<=115;
				end
			end
			5604: begin
				if(in == 0) begin
					state<=5615;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=1726;
					out<=118;
				end
				if(in == 3) begin
					state<=7516;
					out<=119;
				end
				if(in == 4) begin
					state<=3627;
					out<=120;
				end
			end
			5605: begin
				if(in == 0) begin
					state<=5616;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=1727;
					out<=123;
				end
				if(in == 3) begin
					state<=7517;
					out<=124;
				end
				if(in == 4) begin
					state<=3628;
					out<=125;
				end
			end
			5606: begin
				if(in == 0) begin
					state<=5607;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=1718;
					out<=128;
				end
				if(in == 3) begin
					state<=7508;
					out<=129;
				end
				if(in == 4) begin
					state<=3619;
					out<=130;
				end
			end
			5607: begin
				if(in == 0) begin
					state<=5618;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=1729;
					out<=133;
				end
				if(in == 3) begin
					state<=7519;
					out<=134;
				end
				if(in == 4) begin
					state<=3630;
					out<=135;
				end
			end
			5608: begin
				if(in == 0) begin
					state<=5619;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=1730;
					out<=138;
				end
				if(in == 3) begin
					state<=7520;
					out<=139;
				end
				if(in == 4) begin
					state<=3631;
					out<=140;
				end
			end
			5609: begin
				if(in == 0) begin
					state<=5620;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=1731;
					out<=143;
				end
				if(in == 3) begin
					state<=7521;
					out<=144;
				end
				if(in == 4) begin
					state<=3632;
					out<=145;
				end
			end
			5610: begin
				if(in == 0) begin
					state<=5621;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=1732;
					out<=148;
				end
				if(in == 3) begin
					state<=7522;
					out<=149;
				end
				if(in == 4) begin
					state<=3633;
					out<=150;
				end
			end
			5611: begin
				if(in == 0) begin
					state<=5622;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=1733;
					out<=153;
				end
				if(in == 3) begin
					state<=7523;
					out<=154;
				end
				if(in == 4) begin
					state<=3634;
					out<=155;
				end
			end
			5612: begin
				if(in == 0) begin
					state<=5623;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=1734;
					out<=158;
				end
				if(in == 3) begin
					state<=7524;
					out<=159;
				end
				if(in == 4) begin
					state<=3635;
					out<=160;
				end
			end
			5613: begin
				if(in == 0) begin
					state<=5624;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=1735;
					out<=163;
				end
				if(in == 3) begin
					state<=7525;
					out<=164;
				end
				if(in == 4) begin
					state<=3636;
					out<=165;
				end
			end
			5614: begin
				if(in == 0) begin
					state<=5625;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=1736;
					out<=168;
				end
				if(in == 3) begin
					state<=7526;
					out<=169;
				end
				if(in == 4) begin
					state<=3637;
					out<=170;
				end
			end
			5615: begin
				if(in == 0) begin
					state<=5626;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=1737;
					out<=173;
				end
				if(in == 3) begin
					state<=7527;
					out<=174;
				end
				if(in == 4) begin
					state<=3638;
					out<=175;
				end
			end
			5616: begin
				if(in == 0) begin
					state<=5617;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=1728;
					out<=178;
				end
				if(in == 3) begin
					state<=7518;
					out<=179;
				end
				if(in == 4) begin
					state<=3629;
					out<=180;
				end
			end
			5617: begin
				if(in == 0) begin
					state<=5628;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=1739;
					out<=183;
				end
				if(in == 3) begin
					state<=7529;
					out<=184;
				end
				if(in == 4) begin
					state<=3640;
					out<=185;
				end
			end
			5618: begin
				if(in == 0) begin
					state<=5629;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=1740;
					out<=188;
				end
				if(in == 3) begin
					state<=7530;
					out<=189;
				end
				if(in == 4) begin
					state<=3641;
					out<=190;
				end
			end
			5619: begin
				if(in == 0) begin
					state<=5630;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=1741;
					out<=193;
				end
				if(in == 3) begin
					state<=7531;
					out<=194;
				end
				if(in == 4) begin
					state<=3642;
					out<=195;
				end
			end
			5620: begin
				if(in == 0) begin
					state<=5631;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=1742;
					out<=198;
				end
				if(in == 3) begin
					state<=7532;
					out<=199;
				end
				if(in == 4) begin
					state<=3643;
					out<=200;
				end
			end
			5621: begin
				if(in == 0) begin
					state<=5632;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=1743;
					out<=203;
				end
				if(in == 3) begin
					state<=7533;
					out<=204;
				end
				if(in == 4) begin
					state<=3644;
					out<=205;
				end
			end
			5622: begin
				if(in == 0) begin
					state<=5633;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=1744;
					out<=208;
				end
				if(in == 3) begin
					state<=7534;
					out<=209;
				end
				if(in == 4) begin
					state<=3645;
					out<=210;
				end
			end
			5623: begin
				if(in == 0) begin
					state<=5634;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=1745;
					out<=213;
				end
				if(in == 3) begin
					state<=7535;
					out<=214;
				end
				if(in == 4) begin
					state<=3646;
					out<=215;
				end
			end
			5624: begin
				if(in == 0) begin
					state<=5635;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=1746;
					out<=218;
				end
				if(in == 3) begin
					state<=7536;
					out<=219;
				end
				if(in == 4) begin
					state<=3647;
					out<=220;
				end
			end
			5625: begin
				if(in == 0) begin
					state<=5636;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=1747;
					out<=223;
				end
				if(in == 3) begin
					state<=7537;
					out<=224;
				end
				if(in == 4) begin
					state<=3648;
					out<=225;
				end
			end
			5626: begin
				if(in == 0) begin
					state<=5627;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=1738;
					out<=228;
				end
				if(in == 3) begin
					state<=7528;
					out<=229;
				end
				if(in == 4) begin
					state<=3639;
					out<=230;
				end
			end
			5627: begin
				if(in == 0) begin
					state<=5638;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=1749;
					out<=233;
				end
				if(in == 3) begin
					state<=7539;
					out<=234;
				end
				if(in == 4) begin
					state<=3650;
					out<=235;
				end
			end
			5628: begin
				if(in == 0) begin
					state<=5639;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=1750;
					out<=238;
				end
				if(in == 3) begin
					state<=7540;
					out<=239;
				end
				if(in == 4) begin
					state<=3651;
					out<=240;
				end
			end
			5629: begin
				if(in == 0) begin
					state<=5640;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=1751;
					out<=243;
				end
				if(in == 3) begin
					state<=7541;
					out<=244;
				end
				if(in == 4) begin
					state<=3652;
					out<=245;
				end
			end
			5630: begin
				if(in == 0) begin
					state<=5641;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=1752;
					out<=248;
				end
				if(in == 3) begin
					state<=7542;
					out<=249;
				end
				if(in == 4) begin
					state<=3653;
					out<=250;
				end
			end
			5631: begin
				if(in == 0) begin
					state<=5642;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=1753;
					out<=253;
				end
				if(in == 3) begin
					state<=7543;
					out<=254;
				end
				if(in == 4) begin
					state<=3654;
					out<=255;
				end
			end
			5632: begin
				if(in == 0) begin
					state<=5643;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=1754;
					out<=2;
				end
				if(in == 3) begin
					state<=7544;
					out<=3;
				end
				if(in == 4) begin
					state<=3655;
					out<=4;
				end
			end
			5633: begin
				if(in == 0) begin
					state<=5644;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=1755;
					out<=7;
				end
				if(in == 3) begin
					state<=7545;
					out<=8;
				end
				if(in == 4) begin
					state<=3656;
					out<=9;
				end
			end
			5634: begin
				if(in == 0) begin
					state<=5645;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=1756;
					out<=12;
				end
				if(in == 3) begin
					state<=7546;
					out<=13;
				end
				if(in == 4) begin
					state<=3657;
					out<=14;
				end
			end
			5635: begin
				if(in == 0) begin
					state<=5646;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=1757;
					out<=17;
				end
				if(in == 3) begin
					state<=7547;
					out<=18;
				end
				if(in == 4) begin
					state<=3658;
					out<=19;
				end
			end
			5636: begin
				if(in == 0) begin
					state<=5637;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=1748;
					out<=22;
				end
				if(in == 3) begin
					state<=7538;
					out<=23;
				end
				if(in == 4) begin
					state<=3649;
					out<=24;
				end
			end
			5637: begin
				if(in == 0) begin
					state<=5648;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=1759;
					out<=27;
				end
				if(in == 3) begin
					state<=7549;
					out<=28;
				end
				if(in == 4) begin
					state<=3660;
					out<=29;
				end
			end
			5638: begin
				if(in == 0) begin
					state<=5649;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=1760;
					out<=32;
				end
				if(in == 3) begin
					state<=7550;
					out<=33;
				end
				if(in == 4) begin
					state<=3661;
					out<=34;
				end
			end
			5639: begin
				if(in == 0) begin
					state<=5650;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=1761;
					out<=37;
				end
				if(in == 3) begin
					state<=7551;
					out<=38;
				end
				if(in == 4) begin
					state<=3662;
					out<=39;
				end
			end
			5640: begin
				if(in == 0) begin
					state<=5651;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=1762;
					out<=42;
				end
				if(in == 3) begin
					state<=7552;
					out<=43;
				end
				if(in == 4) begin
					state<=3663;
					out<=44;
				end
			end
			5641: begin
				if(in == 0) begin
					state<=5652;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=1763;
					out<=47;
				end
				if(in == 3) begin
					state<=7553;
					out<=48;
				end
				if(in == 4) begin
					state<=3664;
					out<=49;
				end
			end
			5642: begin
				if(in == 0) begin
					state<=5653;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=1764;
					out<=52;
				end
				if(in == 3) begin
					state<=7554;
					out<=53;
				end
				if(in == 4) begin
					state<=3665;
					out<=54;
				end
			end
			5643: begin
				if(in == 0) begin
					state<=5654;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=1765;
					out<=57;
				end
				if(in == 3) begin
					state<=7555;
					out<=58;
				end
				if(in == 4) begin
					state<=3666;
					out<=59;
				end
			end
			5644: begin
				if(in == 0) begin
					state<=5655;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=1766;
					out<=62;
				end
				if(in == 3) begin
					state<=7556;
					out<=63;
				end
				if(in == 4) begin
					state<=3667;
					out<=64;
				end
			end
			5645: begin
				if(in == 0) begin
					state<=5656;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=1767;
					out<=67;
				end
				if(in == 3) begin
					state<=7557;
					out<=68;
				end
				if(in == 4) begin
					state<=3668;
					out<=69;
				end
			end
			5646: begin
				if(in == 0) begin
					state<=5647;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=1758;
					out<=72;
				end
				if(in == 3) begin
					state<=7548;
					out<=73;
				end
				if(in == 4) begin
					state<=3659;
					out<=74;
				end
			end
			5647: begin
				if(in == 0) begin
					state<=5658;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=1769;
					out<=77;
				end
				if(in == 3) begin
					state<=7559;
					out<=78;
				end
				if(in == 4) begin
					state<=3670;
					out<=79;
				end
			end
			5648: begin
				if(in == 0) begin
					state<=5659;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=1770;
					out<=82;
				end
				if(in == 3) begin
					state<=7560;
					out<=83;
				end
				if(in == 4) begin
					state<=3671;
					out<=84;
				end
			end
			5649: begin
				if(in == 0) begin
					state<=5660;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=1771;
					out<=87;
				end
				if(in == 3) begin
					state<=7561;
					out<=88;
				end
				if(in == 4) begin
					state<=3672;
					out<=89;
				end
			end
			5650: begin
				if(in == 0) begin
					state<=5661;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=1772;
					out<=92;
				end
				if(in == 3) begin
					state<=7562;
					out<=93;
				end
				if(in == 4) begin
					state<=3673;
					out<=94;
				end
			end
			5651: begin
				if(in == 0) begin
					state<=5662;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=1773;
					out<=97;
				end
				if(in == 3) begin
					state<=7563;
					out<=98;
				end
				if(in == 4) begin
					state<=3674;
					out<=99;
				end
			end
			5652: begin
				if(in == 0) begin
					state<=5663;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=1774;
					out<=102;
				end
				if(in == 3) begin
					state<=7564;
					out<=103;
				end
				if(in == 4) begin
					state<=3675;
					out<=104;
				end
			end
			5653: begin
				if(in == 0) begin
					state<=5664;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=1775;
					out<=107;
				end
				if(in == 3) begin
					state<=7565;
					out<=108;
				end
				if(in == 4) begin
					state<=3676;
					out<=109;
				end
			end
			5654: begin
				if(in == 0) begin
					state<=5665;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=1776;
					out<=112;
				end
				if(in == 3) begin
					state<=7566;
					out<=113;
				end
				if(in == 4) begin
					state<=3677;
					out<=114;
				end
			end
			5655: begin
				if(in == 0) begin
					state<=5666;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=1777;
					out<=117;
				end
				if(in == 3) begin
					state<=7567;
					out<=118;
				end
				if(in == 4) begin
					state<=3678;
					out<=119;
				end
			end
			5656: begin
				if(in == 0) begin
					state<=5657;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=1768;
					out<=122;
				end
				if(in == 3) begin
					state<=7558;
					out<=123;
				end
				if(in == 4) begin
					state<=3669;
					out<=124;
				end
			end
			5657: begin
				if(in == 0) begin
					state<=5668;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=1779;
					out<=127;
				end
				if(in == 3) begin
					state<=7569;
					out<=128;
				end
				if(in == 4) begin
					state<=3680;
					out<=129;
				end
			end
			5658: begin
				if(in == 0) begin
					state<=5669;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=1780;
					out<=132;
				end
				if(in == 3) begin
					state<=7570;
					out<=133;
				end
				if(in == 4) begin
					state<=3681;
					out<=134;
				end
			end
			5659: begin
				if(in == 0) begin
					state<=5670;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=1781;
					out<=137;
				end
				if(in == 3) begin
					state<=7571;
					out<=138;
				end
				if(in == 4) begin
					state<=3682;
					out<=139;
				end
			end
			5660: begin
				if(in == 0) begin
					state<=5671;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=1782;
					out<=142;
				end
				if(in == 3) begin
					state<=7572;
					out<=143;
				end
				if(in == 4) begin
					state<=3683;
					out<=144;
				end
			end
			5661: begin
				if(in == 0) begin
					state<=5672;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=1783;
					out<=147;
				end
				if(in == 3) begin
					state<=7573;
					out<=148;
				end
				if(in == 4) begin
					state<=3684;
					out<=149;
				end
			end
			5662: begin
				if(in == 0) begin
					state<=5673;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=1784;
					out<=152;
				end
				if(in == 3) begin
					state<=7574;
					out<=153;
				end
				if(in == 4) begin
					state<=3685;
					out<=154;
				end
			end
			5663: begin
				if(in == 0) begin
					state<=5674;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=1785;
					out<=157;
				end
				if(in == 3) begin
					state<=7575;
					out<=158;
				end
				if(in == 4) begin
					state<=3686;
					out<=159;
				end
			end
			5664: begin
				if(in == 0) begin
					state<=5675;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=1786;
					out<=162;
				end
				if(in == 3) begin
					state<=7576;
					out<=163;
				end
				if(in == 4) begin
					state<=3687;
					out<=164;
				end
			end
			5665: begin
				if(in == 0) begin
					state<=5676;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=1787;
					out<=167;
				end
				if(in == 3) begin
					state<=7577;
					out<=168;
				end
				if(in == 4) begin
					state<=3688;
					out<=169;
				end
			end
			5666: begin
				if(in == 0) begin
					state<=5667;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=1778;
					out<=172;
				end
				if(in == 3) begin
					state<=7568;
					out<=173;
				end
				if(in == 4) begin
					state<=3679;
					out<=174;
				end
			end
			5667: begin
				if(in == 0) begin
					state<=5678;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=1789;
					out<=177;
				end
				if(in == 3) begin
					state<=7579;
					out<=178;
				end
				if(in == 4) begin
					state<=3690;
					out<=179;
				end
			end
			5668: begin
				if(in == 0) begin
					state<=5679;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=1790;
					out<=182;
				end
				if(in == 3) begin
					state<=7580;
					out<=183;
				end
				if(in == 4) begin
					state<=3691;
					out<=184;
				end
			end
			5669: begin
				if(in == 0) begin
					state<=5680;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=1791;
					out<=187;
				end
				if(in == 3) begin
					state<=7581;
					out<=188;
				end
				if(in == 4) begin
					state<=3692;
					out<=189;
				end
			end
			5670: begin
				if(in == 0) begin
					state<=5681;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=1792;
					out<=192;
				end
				if(in == 3) begin
					state<=7582;
					out<=193;
				end
				if(in == 4) begin
					state<=3693;
					out<=194;
				end
			end
			5671: begin
				if(in == 0) begin
					state<=5682;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=1793;
					out<=197;
				end
				if(in == 3) begin
					state<=7583;
					out<=198;
				end
				if(in == 4) begin
					state<=3694;
					out<=199;
				end
			end
			5672: begin
				if(in == 0) begin
					state<=5683;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=1794;
					out<=202;
				end
				if(in == 3) begin
					state<=7584;
					out<=203;
				end
				if(in == 4) begin
					state<=3695;
					out<=204;
				end
			end
			5673: begin
				if(in == 0) begin
					state<=5684;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=1795;
					out<=207;
				end
				if(in == 3) begin
					state<=7585;
					out<=208;
				end
				if(in == 4) begin
					state<=3696;
					out<=209;
				end
			end
			5674: begin
				if(in == 0) begin
					state<=5685;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=1796;
					out<=212;
				end
				if(in == 3) begin
					state<=7586;
					out<=213;
				end
				if(in == 4) begin
					state<=3697;
					out<=214;
				end
			end
			5675: begin
				if(in == 0) begin
					state<=5686;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=1797;
					out<=217;
				end
				if(in == 3) begin
					state<=7587;
					out<=218;
				end
				if(in == 4) begin
					state<=3698;
					out<=219;
				end
			end
			5676: begin
				if(in == 0) begin
					state<=5677;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=1788;
					out<=222;
				end
				if(in == 3) begin
					state<=7578;
					out<=223;
				end
				if(in == 4) begin
					state<=3689;
					out<=224;
				end
			end
			5677: begin
				if(in == 0) begin
					state<=5688;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=1799;
					out<=227;
				end
				if(in == 3) begin
					state<=7589;
					out<=228;
				end
				if(in == 4) begin
					state<=3700;
					out<=229;
				end
			end
			5678: begin
				if(in == 0) begin
					state<=5689;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=1800;
					out<=232;
				end
				if(in == 3) begin
					state<=7590;
					out<=233;
				end
				if(in == 4) begin
					state<=3701;
					out<=234;
				end
			end
			5679: begin
				if(in == 0) begin
					state<=5690;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=1801;
					out<=237;
				end
				if(in == 3) begin
					state<=7591;
					out<=238;
				end
				if(in == 4) begin
					state<=3702;
					out<=239;
				end
			end
			5680: begin
				if(in == 0) begin
					state<=5691;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=1802;
					out<=242;
				end
				if(in == 3) begin
					state<=7592;
					out<=243;
				end
				if(in == 4) begin
					state<=3703;
					out<=244;
				end
			end
			5681: begin
				if(in == 0) begin
					state<=5692;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=1803;
					out<=247;
				end
				if(in == 3) begin
					state<=7593;
					out<=248;
				end
				if(in == 4) begin
					state<=3704;
					out<=249;
				end
			end
			5682: begin
				if(in == 0) begin
					state<=5693;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=1804;
					out<=252;
				end
				if(in == 3) begin
					state<=7594;
					out<=253;
				end
				if(in == 4) begin
					state<=3705;
					out<=254;
				end
			end
			5683: begin
				if(in == 0) begin
					state<=5694;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=1805;
					out<=1;
				end
				if(in == 3) begin
					state<=7595;
					out<=2;
				end
				if(in == 4) begin
					state<=3706;
					out<=3;
				end
			end
			5684: begin
				if(in == 0) begin
					state<=5695;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=1806;
					out<=6;
				end
				if(in == 3) begin
					state<=7596;
					out<=7;
				end
				if(in == 4) begin
					state<=3707;
					out<=8;
				end
			end
			5685: begin
				if(in == 0) begin
					state<=5696;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=1807;
					out<=11;
				end
				if(in == 3) begin
					state<=7597;
					out<=12;
				end
				if(in == 4) begin
					state<=3708;
					out<=13;
				end
			end
			5686: begin
				if(in == 0) begin
					state<=5687;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=1798;
					out<=16;
				end
				if(in == 3) begin
					state<=7588;
					out<=17;
				end
				if(in == 4) begin
					state<=3699;
					out<=18;
				end
			end
			5687: begin
				if(in == 0) begin
					state<=5698;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=1809;
					out<=21;
				end
				if(in == 3) begin
					state<=7599;
					out<=22;
				end
				if(in == 4) begin
					state<=3710;
					out<=23;
				end
			end
			5688: begin
				if(in == 0) begin
					state<=5699;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=1810;
					out<=26;
				end
				if(in == 3) begin
					state<=7600;
					out<=27;
				end
				if(in == 4) begin
					state<=3711;
					out<=28;
				end
			end
			5689: begin
				if(in == 0) begin
					state<=5700;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=1811;
					out<=31;
				end
				if(in == 3) begin
					state<=7601;
					out<=32;
				end
				if(in == 4) begin
					state<=3712;
					out<=33;
				end
			end
			5690: begin
				if(in == 0) begin
					state<=5701;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=1812;
					out<=36;
				end
				if(in == 3) begin
					state<=7602;
					out<=37;
				end
				if(in == 4) begin
					state<=3713;
					out<=38;
				end
			end
			5691: begin
				if(in == 0) begin
					state<=5702;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=1813;
					out<=41;
				end
				if(in == 3) begin
					state<=7603;
					out<=42;
				end
				if(in == 4) begin
					state<=3714;
					out<=43;
				end
			end
			5692: begin
				if(in == 0) begin
					state<=5703;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=1814;
					out<=46;
				end
				if(in == 3) begin
					state<=7604;
					out<=47;
				end
				if(in == 4) begin
					state<=3715;
					out<=48;
				end
			end
			5693: begin
				if(in == 0) begin
					state<=5704;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=1815;
					out<=51;
				end
				if(in == 3) begin
					state<=7605;
					out<=52;
				end
				if(in == 4) begin
					state<=3716;
					out<=53;
				end
			end
			5694: begin
				if(in == 0) begin
					state<=5705;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=1816;
					out<=56;
				end
				if(in == 3) begin
					state<=7606;
					out<=57;
				end
				if(in == 4) begin
					state<=3717;
					out<=58;
				end
			end
			5695: begin
				if(in == 0) begin
					state<=5706;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=1817;
					out<=61;
				end
				if(in == 3) begin
					state<=7607;
					out<=62;
				end
				if(in == 4) begin
					state<=3718;
					out<=63;
				end
			end
			5696: begin
				if(in == 0) begin
					state<=5697;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=1808;
					out<=66;
				end
				if(in == 3) begin
					state<=7598;
					out<=67;
				end
				if(in == 4) begin
					state<=3709;
					out<=68;
				end
			end
			5697: begin
				if(in == 0) begin
					state<=5708;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=1819;
					out<=71;
				end
				if(in == 3) begin
					state<=7609;
					out<=72;
				end
				if(in == 4) begin
					state<=3720;
					out<=73;
				end
			end
			5698: begin
				if(in == 0) begin
					state<=5709;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=1820;
					out<=76;
				end
				if(in == 3) begin
					state<=7610;
					out<=77;
				end
				if(in == 4) begin
					state<=3721;
					out<=78;
				end
			end
			5699: begin
				if(in == 0) begin
					state<=5710;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=1821;
					out<=81;
				end
				if(in == 3) begin
					state<=7611;
					out<=82;
				end
				if(in == 4) begin
					state<=3722;
					out<=83;
				end
			end
			5700: begin
				if(in == 0) begin
					state<=5711;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=1822;
					out<=86;
				end
				if(in == 3) begin
					state<=7612;
					out<=87;
				end
				if(in == 4) begin
					state<=3723;
					out<=88;
				end
			end
			5701: begin
				if(in == 0) begin
					state<=5712;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=1823;
					out<=91;
				end
				if(in == 3) begin
					state<=7613;
					out<=92;
				end
				if(in == 4) begin
					state<=3724;
					out<=93;
				end
			end
			5702: begin
				if(in == 0) begin
					state<=5713;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=1824;
					out<=96;
				end
				if(in == 3) begin
					state<=7614;
					out<=97;
				end
				if(in == 4) begin
					state<=3725;
					out<=98;
				end
			end
			5703: begin
				if(in == 0) begin
					state<=5714;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=1825;
					out<=101;
				end
				if(in == 3) begin
					state<=7615;
					out<=102;
				end
				if(in == 4) begin
					state<=3726;
					out<=103;
				end
			end
			5704: begin
				if(in == 0) begin
					state<=5715;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=1826;
					out<=106;
				end
				if(in == 3) begin
					state<=7616;
					out<=107;
				end
				if(in == 4) begin
					state<=3727;
					out<=108;
				end
			end
			5705: begin
				if(in == 0) begin
					state<=5716;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=1827;
					out<=111;
				end
				if(in == 3) begin
					state<=7617;
					out<=112;
				end
				if(in == 4) begin
					state<=3728;
					out<=113;
				end
			end
			5706: begin
				if(in == 0) begin
					state<=5707;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=1818;
					out<=116;
				end
				if(in == 3) begin
					state<=7608;
					out<=117;
				end
				if(in == 4) begin
					state<=3719;
					out<=118;
				end
			end
			5707: begin
				if(in == 0) begin
					state<=5718;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=1829;
					out<=121;
				end
				if(in == 3) begin
					state<=7619;
					out<=122;
				end
				if(in == 4) begin
					state<=3730;
					out<=123;
				end
			end
			5708: begin
				if(in == 0) begin
					state<=5719;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=1830;
					out<=126;
				end
				if(in == 3) begin
					state<=7620;
					out<=127;
				end
				if(in == 4) begin
					state<=3731;
					out<=128;
				end
			end
			5709: begin
				if(in == 0) begin
					state<=5720;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=1831;
					out<=131;
				end
				if(in == 3) begin
					state<=7621;
					out<=132;
				end
				if(in == 4) begin
					state<=3732;
					out<=133;
				end
			end
			5710: begin
				if(in == 0) begin
					state<=5721;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=1832;
					out<=136;
				end
				if(in == 3) begin
					state<=7622;
					out<=137;
				end
				if(in == 4) begin
					state<=3733;
					out<=138;
				end
			end
			5711: begin
				if(in == 0) begin
					state<=5722;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=1833;
					out<=141;
				end
				if(in == 3) begin
					state<=7623;
					out<=142;
				end
				if(in == 4) begin
					state<=3734;
					out<=143;
				end
			end
			5712: begin
				if(in == 0) begin
					state<=5723;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=1834;
					out<=146;
				end
				if(in == 3) begin
					state<=7624;
					out<=147;
				end
				if(in == 4) begin
					state<=3735;
					out<=148;
				end
			end
			5713: begin
				if(in == 0) begin
					state<=5724;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=1835;
					out<=151;
				end
				if(in == 3) begin
					state<=7625;
					out<=152;
				end
				if(in == 4) begin
					state<=3736;
					out<=153;
				end
			end
			5714: begin
				if(in == 0) begin
					state<=5725;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=1836;
					out<=156;
				end
				if(in == 3) begin
					state<=7626;
					out<=157;
				end
				if(in == 4) begin
					state<=3737;
					out<=158;
				end
			end
			5715: begin
				if(in == 0) begin
					state<=5726;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=1837;
					out<=161;
				end
				if(in == 3) begin
					state<=7627;
					out<=162;
				end
				if(in == 4) begin
					state<=3738;
					out<=163;
				end
			end
			5716: begin
				if(in == 0) begin
					state<=5717;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=1828;
					out<=166;
				end
				if(in == 3) begin
					state<=7618;
					out<=167;
				end
				if(in == 4) begin
					state<=3729;
					out<=168;
				end
			end
			5717: begin
				if(in == 0) begin
					state<=5728;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=1839;
					out<=171;
				end
				if(in == 3) begin
					state<=7629;
					out<=172;
				end
				if(in == 4) begin
					state<=3740;
					out<=173;
				end
			end
			5718: begin
				if(in == 0) begin
					state<=5729;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=1840;
					out<=176;
				end
				if(in == 3) begin
					state<=7630;
					out<=177;
				end
				if(in == 4) begin
					state<=3741;
					out<=178;
				end
			end
			5719: begin
				if(in == 0) begin
					state<=5730;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=1841;
					out<=181;
				end
				if(in == 3) begin
					state<=7631;
					out<=182;
				end
				if(in == 4) begin
					state<=3742;
					out<=183;
				end
			end
			5720: begin
				if(in == 0) begin
					state<=5731;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=1842;
					out<=186;
				end
				if(in == 3) begin
					state<=7632;
					out<=187;
				end
				if(in == 4) begin
					state<=3743;
					out<=188;
				end
			end
			5721: begin
				if(in == 0) begin
					state<=5732;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=1843;
					out<=191;
				end
				if(in == 3) begin
					state<=7633;
					out<=192;
				end
				if(in == 4) begin
					state<=3744;
					out<=193;
				end
			end
			5722: begin
				if(in == 0) begin
					state<=5733;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=1844;
					out<=196;
				end
				if(in == 3) begin
					state<=7634;
					out<=197;
				end
				if(in == 4) begin
					state<=3745;
					out<=198;
				end
			end
			5723: begin
				if(in == 0) begin
					state<=5734;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=1845;
					out<=201;
				end
				if(in == 3) begin
					state<=7635;
					out<=202;
				end
				if(in == 4) begin
					state<=3746;
					out<=203;
				end
			end
			5724: begin
				if(in == 0) begin
					state<=5735;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=1846;
					out<=206;
				end
				if(in == 3) begin
					state<=7636;
					out<=207;
				end
				if(in == 4) begin
					state<=3747;
					out<=208;
				end
			end
			5725: begin
				if(in == 0) begin
					state<=5736;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=1847;
					out<=211;
				end
				if(in == 3) begin
					state<=7637;
					out<=212;
				end
				if(in == 4) begin
					state<=3748;
					out<=213;
				end
			end
			5726: begin
				if(in == 0) begin
					state<=5727;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=1838;
					out<=216;
				end
				if(in == 3) begin
					state<=7628;
					out<=217;
				end
				if(in == 4) begin
					state<=3739;
					out<=218;
				end
			end
			5727: begin
				if(in == 0) begin
					state<=5738;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=1849;
					out<=221;
				end
				if(in == 3) begin
					state<=7639;
					out<=222;
				end
				if(in == 4) begin
					state<=3750;
					out<=223;
				end
			end
			5728: begin
				if(in == 0) begin
					state<=5739;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=1850;
					out<=226;
				end
				if(in == 3) begin
					state<=7640;
					out<=227;
				end
				if(in == 4) begin
					state<=3751;
					out<=228;
				end
			end
			5729: begin
				if(in == 0) begin
					state<=5740;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=1851;
					out<=231;
				end
				if(in == 3) begin
					state<=7641;
					out<=232;
				end
				if(in == 4) begin
					state<=3752;
					out<=233;
				end
			end
			5730: begin
				if(in == 0) begin
					state<=5741;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=1852;
					out<=236;
				end
				if(in == 3) begin
					state<=7642;
					out<=237;
				end
				if(in == 4) begin
					state<=3753;
					out<=238;
				end
			end
			5731: begin
				if(in == 0) begin
					state<=5742;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=1853;
					out<=241;
				end
				if(in == 3) begin
					state<=7643;
					out<=242;
				end
				if(in == 4) begin
					state<=3754;
					out<=243;
				end
			end
			5732: begin
				if(in == 0) begin
					state<=5743;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=1854;
					out<=246;
				end
				if(in == 3) begin
					state<=7644;
					out<=247;
				end
				if(in == 4) begin
					state<=3755;
					out<=248;
				end
			end
			5733: begin
				if(in == 0) begin
					state<=5744;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=1855;
					out<=251;
				end
				if(in == 3) begin
					state<=7645;
					out<=252;
				end
				if(in == 4) begin
					state<=3756;
					out<=253;
				end
			end
			5734: begin
				if(in == 0) begin
					state<=5745;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=1856;
					out<=0;
				end
				if(in == 3) begin
					state<=7646;
					out<=1;
				end
				if(in == 4) begin
					state<=3757;
					out<=2;
				end
			end
			5735: begin
				if(in == 0) begin
					state<=5746;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=1857;
					out<=5;
				end
				if(in == 3) begin
					state<=7647;
					out<=6;
				end
				if(in == 4) begin
					state<=3758;
					out<=7;
				end
			end
			5736: begin
				if(in == 0) begin
					state<=5737;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=1848;
					out<=10;
				end
				if(in == 3) begin
					state<=7638;
					out<=11;
				end
				if(in == 4) begin
					state<=3749;
					out<=12;
				end
			end
			5737: begin
				if(in == 0) begin
					state<=5748;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=1859;
					out<=15;
				end
				if(in == 3) begin
					state<=7649;
					out<=16;
				end
				if(in == 4) begin
					state<=3760;
					out<=17;
				end
			end
			5738: begin
				if(in == 0) begin
					state<=5749;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=1860;
					out<=20;
				end
				if(in == 3) begin
					state<=7650;
					out<=21;
				end
				if(in == 4) begin
					state<=3761;
					out<=22;
				end
			end
			5739: begin
				if(in == 0) begin
					state<=5750;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=1861;
					out<=25;
				end
				if(in == 3) begin
					state<=7651;
					out<=26;
				end
				if(in == 4) begin
					state<=3762;
					out<=27;
				end
			end
			5740: begin
				if(in == 0) begin
					state<=5751;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=1862;
					out<=30;
				end
				if(in == 3) begin
					state<=7652;
					out<=31;
				end
				if(in == 4) begin
					state<=3763;
					out<=32;
				end
			end
			5741: begin
				if(in == 0) begin
					state<=5752;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=1863;
					out<=35;
				end
				if(in == 3) begin
					state<=7653;
					out<=36;
				end
				if(in == 4) begin
					state<=3764;
					out<=37;
				end
			end
			5742: begin
				if(in == 0) begin
					state<=5753;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=1864;
					out<=40;
				end
				if(in == 3) begin
					state<=7654;
					out<=41;
				end
				if(in == 4) begin
					state<=3765;
					out<=42;
				end
			end
			5743: begin
				if(in == 0) begin
					state<=5754;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=1865;
					out<=45;
				end
				if(in == 3) begin
					state<=7655;
					out<=46;
				end
				if(in == 4) begin
					state<=3766;
					out<=47;
				end
			end
			5744: begin
				if(in == 0) begin
					state<=5755;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=1866;
					out<=50;
				end
				if(in == 3) begin
					state<=7656;
					out<=51;
				end
				if(in == 4) begin
					state<=3767;
					out<=52;
				end
			end
			5745: begin
				if(in == 0) begin
					state<=5756;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=1867;
					out<=55;
				end
				if(in == 3) begin
					state<=7657;
					out<=56;
				end
				if(in == 4) begin
					state<=3768;
					out<=57;
				end
			end
			5746: begin
				if(in == 0) begin
					state<=5747;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=1858;
					out<=60;
				end
				if(in == 3) begin
					state<=7648;
					out<=61;
				end
				if(in == 4) begin
					state<=3759;
					out<=62;
				end
			end
			5747: begin
				if(in == 0) begin
					state<=5758;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=1869;
					out<=65;
				end
				if(in == 3) begin
					state<=7659;
					out<=66;
				end
				if(in == 4) begin
					state<=3770;
					out<=67;
				end
			end
			5748: begin
				if(in == 0) begin
					state<=5759;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=1870;
					out<=70;
				end
				if(in == 3) begin
					state<=7660;
					out<=71;
				end
				if(in == 4) begin
					state<=3771;
					out<=72;
				end
			end
			5749: begin
				if(in == 0) begin
					state<=5760;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=1871;
					out<=75;
				end
				if(in == 3) begin
					state<=7661;
					out<=76;
				end
				if(in == 4) begin
					state<=3772;
					out<=77;
				end
			end
			5750: begin
				if(in == 0) begin
					state<=5761;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=1872;
					out<=80;
				end
				if(in == 3) begin
					state<=7662;
					out<=81;
				end
				if(in == 4) begin
					state<=3773;
					out<=82;
				end
			end
			5751: begin
				if(in == 0) begin
					state<=5762;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=1873;
					out<=85;
				end
				if(in == 3) begin
					state<=7663;
					out<=86;
				end
				if(in == 4) begin
					state<=3774;
					out<=87;
				end
			end
			5752: begin
				if(in == 0) begin
					state<=5763;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=1874;
					out<=90;
				end
				if(in == 3) begin
					state<=7664;
					out<=91;
				end
				if(in == 4) begin
					state<=3775;
					out<=92;
				end
			end
			5753: begin
				if(in == 0) begin
					state<=5764;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=1875;
					out<=95;
				end
				if(in == 3) begin
					state<=7665;
					out<=96;
				end
				if(in == 4) begin
					state<=3776;
					out<=97;
				end
			end
			5754: begin
				if(in == 0) begin
					state<=5765;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=1876;
					out<=100;
				end
				if(in == 3) begin
					state<=7666;
					out<=101;
				end
				if(in == 4) begin
					state<=3777;
					out<=102;
				end
			end
			5755: begin
				if(in == 0) begin
					state<=5766;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=1877;
					out<=105;
				end
				if(in == 3) begin
					state<=7667;
					out<=106;
				end
				if(in == 4) begin
					state<=3778;
					out<=107;
				end
			end
			5756: begin
				if(in == 0) begin
					state<=5757;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=1868;
					out<=110;
				end
				if(in == 3) begin
					state<=7658;
					out<=111;
				end
				if(in == 4) begin
					state<=3769;
					out<=112;
				end
			end
			5757: begin
				if(in == 0) begin
					state<=5768;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=1879;
					out<=115;
				end
				if(in == 3) begin
					state<=7669;
					out<=116;
				end
				if(in == 4) begin
					state<=3780;
					out<=117;
				end
			end
			5758: begin
				if(in == 0) begin
					state<=5769;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=1880;
					out<=120;
				end
				if(in == 3) begin
					state<=7670;
					out<=121;
				end
				if(in == 4) begin
					state<=3781;
					out<=122;
				end
			end
			5759: begin
				if(in == 0) begin
					state<=5770;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=1881;
					out<=125;
				end
				if(in == 3) begin
					state<=7671;
					out<=126;
				end
				if(in == 4) begin
					state<=3782;
					out<=127;
				end
			end
			5760: begin
				if(in == 0) begin
					state<=5771;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=1882;
					out<=130;
				end
				if(in == 3) begin
					state<=7672;
					out<=131;
				end
				if(in == 4) begin
					state<=3783;
					out<=132;
				end
			end
			5761: begin
				if(in == 0) begin
					state<=5772;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=1883;
					out<=135;
				end
				if(in == 3) begin
					state<=7673;
					out<=136;
				end
				if(in == 4) begin
					state<=3784;
					out<=137;
				end
			end
			5762: begin
				if(in == 0) begin
					state<=5773;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=1884;
					out<=140;
				end
				if(in == 3) begin
					state<=7674;
					out<=141;
				end
				if(in == 4) begin
					state<=3785;
					out<=142;
				end
			end
			5763: begin
				if(in == 0) begin
					state<=5774;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=1885;
					out<=145;
				end
				if(in == 3) begin
					state<=7675;
					out<=146;
				end
				if(in == 4) begin
					state<=3786;
					out<=147;
				end
			end
			5764: begin
				if(in == 0) begin
					state<=5775;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=1886;
					out<=150;
				end
				if(in == 3) begin
					state<=7676;
					out<=151;
				end
				if(in == 4) begin
					state<=3787;
					out<=152;
				end
			end
			5765: begin
				if(in == 0) begin
					state<=5776;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=1887;
					out<=155;
				end
				if(in == 3) begin
					state<=7677;
					out<=156;
				end
				if(in == 4) begin
					state<=3788;
					out<=157;
				end
			end
			5766: begin
				if(in == 0) begin
					state<=5767;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=1878;
					out<=160;
				end
				if(in == 3) begin
					state<=7668;
					out<=161;
				end
				if(in == 4) begin
					state<=3779;
					out<=162;
				end
			end
			5767: begin
				if(in == 0) begin
					state<=5778;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=1889;
					out<=165;
				end
				if(in == 3) begin
					state<=7679;
					out<=166;
				end
				if(in == 4) begin
					state<=3790;
					out<=167;
				end
			end
			5768: begin
				if(in == 0) begin
					state<=5779;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=1890;
					out<=170;
				end
				if(in == 3) begin
					state<=7680;
					out<=171;
				end
				if(in == 4) begin
					state<=3791;
					out<=172;
				end
			end
			5769: begin
				if(in == 0) begin
					state<=5780;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=1891;
					out<=175;
				end
				if(in == 3) begin
					state<=7681;
					out<=176;
				end
				if(in == 4) begin
					state<=3792;
					out<=177;
				end
			end
			5770: begin
				if(in == 0) begin
					state<=5781;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=1892;
					out<=180;
				end
				if(in == 3) begin
					state<=7682;
					out<=181;
				end
				if(in == 4) begin
					state<=3793;
					out<=182;
				end
			end
			5771: begin
				if(in == 0) begin
					state<=5782;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=1893;
					out<=185;
				end
				if(in == 3) begin
					state<=7683;
					out<=186;
				end
				if(in == 4) begin
					state<=3794;
					out<=187;
				end
			end
			5772: begin
				if(in == 0) begin
					state<=5783;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=1894;
					out<=190;
				end
				if(in == 3) begin
					state<=7684;
					out<=191;
				end
				if(in == 4) begin
					state<=3795;
					out<=192;
				end
			end
			5773: begin
				if(in == 0) begin
					state<=5784;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=1895;
					out<=195;
				end
				if(in == 3) begin
					state<=7685;
					out<=196;
				end
				if(in == 4) begin
					state<=3796;
					out<=197;
				end
			end
			5774: begin
				if(in == 0) begin
					state<=5785;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=1896;
					out<=200;
				end
				if(in == 3) begin
					state<=7686;
					out<=201;
				end
				if(in == 4) begin
					state<=3797;
					out<=202;
				end
			end
			5775: begin
				if(in == 0) begin
					state<=5786;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=1897;
					out<=205;
				end
				if(in == 3) begin
					state<=7687;
					out<=206;
				end
				if(in == 4) begin
					state<=3798;
					out<=207;
				end
			end
			5776: begin
				if(in == 0) begin
					state<=5777;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=1888;
					out<=210;
				end
				if(in == 3) begin
					state<=7678;
					out<=211;
				end
				if(in == 4) begin
					state<=3789;
					out<=212;
				end
			end
			5777: begin
				if(in == 0) begin
					state<=5788;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=1899;
					out<=215;
				end
				if(in == 3) begin
					state<=7689;
					out<=216;
				end
				if(in == 4) begin
					state<=3800;
					out<=217;
				end
			end
			5778: begin
				if(in == 0) begin
					state<=5789;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=1900;
					out<=220;
				end
				if(in == 3) begin
					state<=7690;
					out<=221;
				end
				if(in == 4) begin
					state<=3801;
					out<=222;
				end
			end
			5779: begin
				if(in == 0) begin
					state<=5790;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=1901;
					out<=225;
				end
				if(in == 3) begin
					state<=7691;
					out<=226;
				end
				if(in == 4) begin
					state<=3802;
					out<=227;
				end
			end
			5780: begin
				if(in == 0) begin
					state<=5791;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=1902;
					out<=230;
				end
				if(in == 3) begin
					state<=7692;
					out<=231;
				end
				if(in == 4) begin
					state<=3803;
					out<=232;
				end
			end
			5781: begin
				if(in == 0) begin
					state<=5792;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=1903;
					out<=235;
				end
				if(in == 3) begin
					state<=7693;
					out<=236;
				end
				if(in == 4) begin
					state<=3804;
					out<=237;
				end
			end
			5782: begin
				if(in == 0) begin
					state<=5793;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=1904;
					out<=240;
				end
				if(in == 3) begin
					state<=7694;
					out<=241;
				end
				if(in == 4) begin
					state<=3805;
					out<=242;
				end
			end
			5783: begin
				if(in == 0) begin
					state<=5794;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=1905;
					out<=245;
				end
				if(in == 3) begin
					state<=7695;
					out<=246;
				end
				if(in == 4) begin
					state<=3806;
					out<=247;
				end
			end
			5784: begin
				if(in == 0) begin
					state<=5795;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=1906;
					out<=250;
				end
				if(in == 3) begin
					state<=7696;
					out<=251;
				end
				if(in == 4) begin
					state<=3807;
					out<=252;
				end
			end
			5785: begin
				if(in == 0) begin
					state<=5796;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=1907;
					out<=255;
				end
				if(in == 3) begin
					state<=7697;
					out<=0;
				end
				if(in == 4) begin
					state<=3808;
					out<=1;
				end
			end
			5786: begin
				if(in == 0) begin
					state<=5787;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=1898;
					out<=4;
				end
				if(in == 3) begin
					state<=7688;
					out<=5;
				end
				if(in == 4) begin
					state<=3799;
					out<=6;
				end
			end
			5787: begin
				if(in == 0) begin
					state<=5798;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=1909;
					out<=9;
				end
				if(in == 3) begin
					state<=7699;
					out<=10;
				end
				if(in == 4) begin
					state<=3810;
					out<=11;
				end
			end
			5788: begin
				if(in == 0) begin
					state<=5799;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=1910;
					out<=14;
				end
				if(in == 3) begin
					state<=7700;
					out<=15;
				end
				if(in == 4) begin
					state<=3811;
					out<=16;
				end
			end
			5789: begin
				if(in == 0) begin
					state<=5800;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=1911;
					out<=19;
				end
				if(in == 3) begin
					state<=7701;
					out<=20;
				end
				if(in == 4) begin
					state<=3812;
					out<=21;
				end
			end
			5790: begin
				if(in == 0) begin
					state<=5801;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=1912;
					out<=24;
				end
				if(in == 3) begin
					state<=7702;
					out<=25;
				end
				if(in == 4) begin
					state<=3813;
					out<=26;
				end
			end
			5791: begin
				if(in == 0) begin
					state<=5802;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=1913;
					out<=29;
				end
				if(in == 3) begin
					state<=7703;
					out<=30;
				end
				if(in == 4) begin
					state<=3814;
					out<=31;
				end
			end
			5792: begin
				if(in == 0) begin
					state<=5803;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=1914;
					out<=34;
				end
				if(in == 3) begin
					state<=7704;
					out<=35;
				end
				if(in == 4) begin
					state<=3815;
					out<=36;
				end
			end
			5793: begin
				if(in == 0) begin
					state<=5804;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=1915;
					out<=39;
				end
				if(in == 3) begin
					state<=7705;
					out<=40;
				end
				if(in == 4) begin
					state<=3816;
					out<=41;
				end
			end
			5794: begin
				if(in == 0) begin
					state<=5805;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=1916;
					out<=44;
				end
				if(in == 3) begin
					state<=7706;
					out<=45;
				end
				if(in == 4) begin
					state<=3817;
					out<=46;
				end
			end
			5795: begin
				if(in == 0) begin
					state<=5806;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=1917;
					out<=49;
				end
				if(in == 3) begin
					state<=7707;
					out<=50;
				end
				if(in == 4) begin
					state<=3818;
					out<=51;
				end
			end
			5796: begin
				if(in == 0) begin
					state<=5797;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=1908;
					out<=54;
				end
				if(in == 3) begin
					state<=7698;
					out<=55;
				end
				if(in == 4) begin
					state<=3809;
					out<=56;
				end
			end
			5797: begin
				if(in == 0) begin
					state<=5808;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=1919;
					out<=59;
				end
				if(in == 3) begin
					state<=7709;
					out<=60;
				end
				if(in == 4) begin
					state<=3820;
					out<=61;
				end
			end
			5798: begin
				if(in == 0) begin
					state<=5809;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=1920;
					out<=64;
				end
				if(in == 3) begin
					state<=7710;
					out<=65;
				end
				if(in == 4) begin
					state<=3821;
					out<=66;
				end
			end
			5799: begin
				if(in == 0) begin
					state<=5810;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=1921;
					out<=69;
				end
				if(in == 3) begin
					state<=7711;
					out<=70;
				end
				if(in == 4) begin
					state<=3822;
					out<=71;
				end
			end
			5800: begin
				if(in == 0) begin
					state<=5811;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=1922;
					out<=74;
				end
				if(in == 3) begin
					state<=7712;
					out<=75;
				end
				if(in == 4) begin
					state<=3823;
					out<=76;
				end
			end
			5801: begin
				if(in == 0) begin
					state<=5812;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=1923;
					out<=79;
				end
				if(in == 3) begin
					state<=7713;
					out<=80;
				end
				if(in == 4) begin
					state<=3824;
					out<=81;
				end
			end
			5802: begin
				if(in == 0) begin
					state<=5813;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=1924;
					out<=84;
				end
				if(in == 3) begin
					state<=7714;
					out<=85;
				end
				if(in == 4) begin
					state<=3825;
					out<=86;
				end
			end
			5803: begin
				if(in == 0) begin
					state<=5814;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=1925;
					out<=89;
				end
				if(in == 3) begin
					state<=7715;
					out<=90;
				end
				if(in == 4) begin
					state<=3826;
					out<=91;
				end
			end
			5804: begin
				if(in == 0) begin
					state<=5815;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=1926;
					out<=94;
				end
				if(in == 3) begin
					state<=7716;
					out<=95;
				end
				if(in == 4) begin
					state<=3827;
					out<=96;
				end
			end
			5805: begin
				if(in == 0) begin
					state<=5816;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=1927;
					out<=99;
				end
				if(in == 3) begin
					state<=7717;
					out<=100;
				end
				if(in == 4) begin
					state<=3828;
					out<=101;
				end
			end
			5806: begin
				if(in == 0) begin
					state<=5807;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=1918;
					out<=104;
				end
				if(in == 3) begin
					state<=7708;
					out<=105;
				end
				if(in == 4) begin
					state<=3819;
					out<=106;
				end
			end
			5807: begin
				if(in == 0) begin
					state<=5818;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=1929;
					out<=109;
				end
				if(in == 3) begin
					state<=7719;
					out<=110;
				end
				if(in == 4) begin
					state<=3830;
					out<=111;
				end
			end
			5808: begin
				if(in == 0) begin
					state<=5819;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=1930;
					out<=114;
				end
				if(in == 3) begin
					state<=7720;
					out<=115;
				end
				if(in == 4) begin
					state<=3831;
					out<=116;
				end
			end
			5809: begin
				if(in == 0) begin
					state<=5820;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=1931;
					out<=119;
				end
				if(in == 3) begin
					state<=7721;
					out<=120;
				end
				if(in == 4) begin
					state<=3832;
					out<=121;
				end
			end
			5810: begin
				if(in == 0) begin
					state<=5821;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=1932;
					out<=124;
				end
				if(in == 3) begin
					state<=7722;
					out<=125;
				end
				if(in == 4) begin
					state<=3833;
					out<=126;
				end
			end
			5811: begin
				if(in == 0) begin
					state<=5822;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=1933;
					out<=129;
				end
				if(in == 3) begin
					state<=7723;
					out<=130;
				end
				if(in == 4) begin
					state<=3834;
					out<=131;
				end
			end
			5812: begin
				if(in == 0) begin
					state<=5823;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=1934;
					out<=134;
				end
				if(in == 3) begin
					state<=7724;
					out<=135;
				end
				if(in == 4) begin
					state<=3835;
					out<=136;
				end
			end
			5813: begin
				if(in == 0) begin
					state<=5824;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=1935;
					out<=139;
				end
				if(in == 3) begin
					state<=7725;
					out<=140;
				end
				if(in == 4) begin
					state<=3836;
					out<=141;
				end
			end
			5814: begin
				if(in == 0) begin
					state<=5825;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=1936;
					out<=144;
				end
				if(in == 3) begin
					state<=7726;
					out<=145;
				end
				if(in == 4) begin
					state<=3837;
					out<=146;
				end
			end
			5815: begin
				if(in == 0) begin
					state<=5826;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=1937;
					out<=149;
				end
				if(in == 3) begin
					state<=7727;
					out<=150;
				end
				if(in == 4) begin
					state<=3838;
					out<=151;
				end
			end
			5816: begin
				if(in == 0) begin
					state<=5817;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=1928;
					out<=154;
				end
				if(in == 3) begin
					state<=7718;
					out<=155;
				end
				if(in == 4) begin
					state<=3829;
					out<=156;
				end
			end
			5817: begin
				if(in == 0) begin
					state<=5828;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=1939;
					out<=159;
				end
				if(in == 3) begin
					state<=7729;
					out<=160;
				end
				if(in == 4) begin
					state<=3840;
					out<=161;
				end
			end
			5818: begin
				if(in == 0) begin
					state<=5829;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=1940;
					out<=164;
				end
				if(in == 3) begin
					state<=7730;
					out<=165;
				end
				if(in == 4) begin
					state<=3841;
					out<=166;
				end
			end
			5819: begin
				if(in == 0) begin
					state<=5830;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=1941;
					out<=169;
				end
				if(in == 3) begin
					state<=7731;
					out<=170;
				end
				if(in == 4) begin
					state<=3842;
					out<=171;
				end
			end
			5820: begin
				if(in == 0) begin
					state<=5831;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=1942;
					out<=174;
				end
				if(in == 3) begin
					state<=7732;
					out<=175;
				end
				if(in == 4) begin
					state<=3843;
					out<=176;
				end
			end
			5821: begin
				if(in == 0) begin
					state<=5832;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=1943;
					out<=179;
				end
				if(in == 3) begin
					state<=7733;
					out<=180;
				end
				if(in == 4) begin
					state<=3844;
					out<=181;
				end
			end
			5822: begin
				if(in == 0) begin
					state<=5833;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=1944;
					out<=184;
				end
				if(in == 3) begin
					state<=7734;
					out<=185;
				end
				if(in == 4) begin
					state<=3845;
					out<=186;
				end
			end
			5823: begin
				if(in == 0) begin
					state<=5834;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=1945;
					out<=189;
				end
				if(in == 3) begin
					state<=7735;
					out<=190;
				end
				if(in == 4) begin
					state<=3846;
					out<=191;
				end
			end
			5824: begin
				if(in == 0) begin
					state<=5835;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=1946;
					out<=194;
				end
				if(in == 3) begin
					state<=7736;
					out<=195;
				end
				if(in == 4) begin
					state<=3847;
					out<=196;
				end
			end
			5825: begin
				if(in == 0) begin
					state<=5836;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=1947;
					out<=199;
				end
				if(in == 3) begin
					state<=7737;
					out<=200;
				end
				if(in == 4) begin
					state<=3848;
					out<=201;
				end
			end
			5826: begin
				if(in == 0) begin
					state<=5827;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=1938;
					out<=204;
				end
				if(in == 3) begin
					state<=7728;
					out<=205;
				end
				if(in == 4) begin
					state<=3839;
					out<=206;
				end
			end
			5827: begin
				if(in == 0) begin
					state<=5838;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=1949;
					out<=209;
				end
				if(in == 3) begin
					state<=7739;
					out<=210;
				end
				if(in == 4) begin
					state<=3850;
					out<=211;
				end
			end
			5828: begin
				if(in == 0) begin
					state<=5839;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=1950;
					out<=214;
				end
				if(in == 3) begin
					state<=7740;
					out<=215;
				end
				if(in == 4) begin
					state<=3851;
					out<=216;
				end
			end
			5829: begin
				if(in == 0) begin
					state<=5840;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=1951;
					out<=219;
				end
				if(in == 3) begin
					state<=7741;
					out<=220;
				end
				if(in == 4) begin
					state<=3852;
					out<=221;
				end
			end
			5830: begin
				if(in == 0) begin
					state<=5841;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=1952;
					out<=224;
				end
				if(in == 3) begin
					state<=7742;
					out<=225;
				end
				if(in == 4) begin
					state<=3853;
					out<=226;
				end
			end
			5831: begin
				if(in == 0) begin
					state<=5842;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=1953;
					out<=229;
				end
				if(in == 3) begin
					state<=7743;
					out<=230;
				end
				if(in == 4) begin
					state<=3854;
					out<=231;
				end
			end
			5832: begin
				if(in == 0) begin
					state<=5843;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=1954;
					out<=234;
				end
				if(in == 3) begin
					state<=7744;
					out<=235;
				end
				if(in == 4) begin
					state<=3855;
					out<=236;
				end
			end
			5833: begin
				if(in == 0) begin
					state<=5844;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=1955;
					out<=239;
				end
				if(in == 3) begin
					state<=7745;
					out<=240;
				end
				if(in == 4) begin
					state<=3856;
					out<=241;
				end
			end
			5834: begin
				if(in == 0) begin
					state<=5845;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=1956;
					out<=244;
				end
				if(in == 3) begin
					state<=7746;
					out<=245;
				end
				if(in == 4) begin
					state<=3857;
					out<=246;
				end
			end
			5835: begin
				if(in == 0) begin
					state<=5846;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=1957;
					out<=249;
				end
				if(in == 3) begin
					state<=7747;
					out<=250;
				end
				if(in == 4) begin
					state<=3858;
					out<=251;
				end
			end
			5836: begin
				if(in == 0) begin
					state<=5837;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=1948;
					out<=254;
				end
				if(in == 3) begin
					state<=7738;
					out<=255;
				end
				if(in == 4) begin
					state<=3849;
					out<=0;
				end
			end
			5837: begin
				if(in == 0) begin
					state<=5848;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=1959;
					out<=3;
				end
				if(in == 3) begin
					state<=7749;
					out<=4;
				end
				if(in == 4) begin
					state<=3860;
					out<=5;
				end
			end
			5838: begin
				if(in == 0) begin
					state<=5849;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=1960;
					out<=8;
				end
				if(in == 3) begin
					state<=7750;
					out<=9;
				end
				if(in == 4) begin
					state<=3861;
					out<=10;
				end
			end
			5839: begin
				if(in == 0) begin
					state<=5850;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=1961;
					out<=13;
				end
				if(in == 3) begin
					state<=7751;
					out<=14;
				end
				if(in == 4) begin
					state<=3862;
					out<=15;
				end
			end
			5840: begin
				if(in == 0) begin
					state<=5851;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=1962;
					out<=18;
				end
				if(in == 3) begin
					state<=7752;
					out<=19;
				end
				if(in == 4) begin
					state<=3863;
					out<=20;
				end
			end
			5841: begin
				if(in == 0) begin
					state<=5852;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=1963;
					out<=23;
				end
				if(in == 3) begin
					state<=7753;
					out<=24;
				end
				if(in == 4) begin
					state<=3864;
					out<=25;
				end
			end
			5842: begin
				if(in == 0) begin
					state<=5853;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=1964;
					out<=28;
				end
				if(in == 3) begin
					state<=7754;
					out<=29;
				end
				if(in == 4) begin
					state<=3865;
					out<=30;
				end
			end
			5843: begin
				if(in == 0) begin
					state<=5854;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=1965;
					out<=33;
				end
				if(in == 3) begin
					state<=7755;
					out<=34;
				end
				if(in == 4) begin
					state<=3866;
					out<=35;
				end
			end
			5844: begin
				if(in == 0) begin
					state<=5855;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=1966;
					out<=38;
				end
				if(in == 3) begin
					state<=7756;
					out<=39;
				end
				if(in == 4) begin
					state<=3867;
					out<=40;
				end
			end
			5845: begin
				if(in == 0) begin
					state<=5856;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=1967;
					out<=43;
				end
				if(in == 3) begin
					state<=7757;
					out<=44;
				end
				if(in == 4) begin
					state<=3868;
					out<=45;
				end
			end
			5846: begin
				if(in == 0) begin
					state<=5847;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=1958;
					out<=48;
				end
				if(in == 3) begin
					state<=7748;
					out<=49;
				end
				if(in == 4) begin
					state<=3859;
					out<=50;
				end
			end
			5847: begin
				if(in == 0) begin
					state<=5858;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=1969;
					out<=53;
				end
				if(in == 3) begin
					state<=7759;
					out<=54;
				end
				if(in == 4) begin
					state<=3870;
					out<=55;
				end
			end
			5848: begin
				if(in == 0) begin
					state<=5859;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=1970;
					out<=58;
				end
				if(in == 3) begin
					state<=7760;
					out<=59;
				end
				if(in == 4) begin
					state<=3871;
					out<=60;
				end
			end
			5849: begin
				if(in == 0) begin
					state<=5860;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=1971;
					out<=63;
				end
				if(in == 3) begin
					state<=7761;
					out<=64;
				end
				if(in == 4) begin
					state<=3872;
					out<=65;
				end
			end
			5850: begin
				if(in == 0) begin
					state<=5861;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=1972;
					out<=68;
				end
				if(in == 3) begin
					state<=7762;
					out<=69;
				end
				if(in == 4) begin
					state<=3873;
					out<=70;
				end
			end
			5851: begin
				if(in == 0) begin
					state<=5862;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=1973;
					out<=73;
				end
				if(in == 3) begin
					state<=7763;
					out<=74;
				end
				if(in == 4) begin
					state<=3874;
					out<=75;
				end
			end
			5852: begin
				if(in == 0) begin
					state<=5863;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=1974;
					out<=78;
				end
				if(in == 3) begin
					state<=7764;
					out<=79;
				end
				if(in == 4) begin
					state<=3875;
					out<=80;
				end
			end
			5853: begin
				if(in == 0) begin
					state<=5864;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=1975;
					out<=83;
				end
				if(in == 3) begin
					state<=7765;
					out<=84;
				end
				if(in == 4) begin
					state<=3876;
					out<=85;
				end
			end
			5854: begin
				if(in == 0) begin
					state<=5865;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=1976;
					out<=88;
				end
				if(in == 3) begin
					state<=7766;
					out<=89;
				end
				if(in == 4) begin
					state<=3877;
					out<=90;
				end
			end
			5855: begin
				if(in == 0) begin
					state<=5866;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=1977;
					out<=93;
				end
				if(in == 3) begin
					state<=7767;
					out<=94;
				end
				if(in == 4) begin
					state<=3878;
					out<=95;
				end
			end
			5856: begin
				if(in == 0) begin
					state<=5857;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=1968;
					out<=98;
				end
				if(in == 3) begin
					state<=7758;
					out<=99;
				end
				if(in == 4) begin
					state<=3869;
					out<=100;
				end
			end
			5857: begin
				if(in == 0) begin
					state<=5868;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=1979;
					out<=103;
				end
				if(in == 3) begin
					state<=7769;
					out<=104;
				end
				if(in == 4) begin
					state<=3880;
					out<=105;
				end
			end
			5858: begin
				if(in == 0) begin
					state<=5869;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=1980;
					out<=108;
				end
				if(in == 3) begin
					state<=7770;
					out<=109;
				end
				if(in == 4) begin
					state<=3881;
					out<=110;
				end
			end
			5859: begin
				if(in == 0) begin
					state<=5870;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=1981;
					out<=113;
				end
				if(in == 3) begin
					state<=7771;
					out<=114;
				end
				if(in == 4) begin
					state<=3882;
					out<=115;
				end
			end
			5860: begin
				if(in == 0) begin
					state<=5871;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=1982;
					out<=118;
				end
				if(in == 3) begin
					state<=7772;
					out<=119;
				end
				if(in == 4) begin
					state<=3883;
					out<=120;
				end
			end
			5861: begin
				if(in == 0) begin
					state<=5872;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=1983;
					out<=123;
				end
				if(in == 3) begin
					state<=7773;
					out<=124;
				end
				if(in == 4) begin
					state<=3884;
					out<=125;
				end
			end
			5862: begin
				if(in == 0) begin
					state<=5873;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=1984;
					out<=128;
				end
				if(in == 3) begin
					state<=7774;
					out<=129;
				end
				if(in == 4) begin
					state<=3885;
					out<=130;
				end
			end
			5863: begin
				if(in == 0) begin
					state<=5874;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=1985;
					out<=133;
				end
				if(in == 3) begin
					state<=7775;
					out<=134;
				end
				if(in == 4) begin
					state<=3886;
					out<=135;
				end
			end
			5864: begin
				if(in == 0) begin
					state<=5875;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=1986;
					out<=138;
				end
				if(in == 3) begin
					state<=7776;
					out<=139;
				end
				if(in == 4) begin
					state<=3887;
					out<=140;
				end
			end
			5865: begin
				if(in == 0) begin
					state<=5876;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=1987;
					out<=143;
				end
				if(in == 3) begin
					state<=7777;
					out<=144;
				end
				if(in == 4) begin
					state<=3888;
					out<=145;
				end
			end
			5866: begin
				if(in == 0) begin
					state<=5867;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=1978;
					out<=148;
				end
				if(in == 3) begin
					state<=7768;
					out<=149;
				end
				if(in == 4) begin
					state<=3879;
					out<=150;
				end
			end
			5867: begin
				if(in == 0) begin
					state<=5878;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=1989;
					out<=153;
				end
				if(in == 3) begin
					state<=7779;
					out<=154;
				end
				if(in == 4) begin
					state<=3890;
					out<=155;
				end
			end
			5868: begin
				if(in == 0) begin
					state<=5879;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=1990;
					out<=158;
				end
				if(in == 3) begin
					state<=7780;
					out<=159;
				end
				if(in == 4) begin
					state<=3891;
					out<=160;
				end
			end
			5869: begin
				if(in == 0) begin
					state<=5880;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=1991;
					out<=163;
				end
				if(in == 3) begin
					state<=7781;
					out<=164;
				end
				if(in == 4) begin
					state<=3892;
					out<=165;
				end
			end
			5870: begin
				if(in == 0) begin
					state<=5881;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=1992;
					out<=168;
				end
				if(in == 3) begin
					state<=7782;
					out<=169;
				end
				if(in == 4) begin
					state<=3893;
					out<=170;
				end
			end
			5871: begin
				if(in == 0) begin
					state<=5882;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=1993;
					out<=173;
				end
				if(in == 3) begin
					state<=7783;
					out<=174;
				end
				if(in == 4) begin
					state<=3894;
					out<=175;
				end
			end
			5872: begin
				if(in == 0) begin
					state<=5883;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=1994;
					out<=178;
				end
				if(in == 3) begin
					state<=7784;
					out<=179;
				end
				if(in == 4) begin
					state<=3895;
					out<=180;
				end
			end
			5873: begin
				if(in == 0) begin
					state<=5884;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=1995;
					out<=183;
				end
				if(in == 3) begin
					state<=7785;
					out<=184;
				end
				if(in == 4) begin
					state<=3896;
					out<=185;
				end
			end
			5874: begin
				if(in == 0) begin
					state<=5885;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=1996;
					out<=188;
				end
				if(in == 3) begin
					state<=7786;
					out<=189;
				end
				if(in == 4) begin
					state<=3897;
					out<=190;
				end
			end
			5875: begin
				if(in == 0) begin
					state<=5886;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=1997;
					out<=193;
				end
				if(in == 3) begin
					state<=7787;
					out<=194;
				end
				if(in == 4) begin
					state<=3898;
					out<=195;
				end
			end
			5876: begin
				if(in == 0) begin
					state<=5877;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=1988;
					out<=198;
				end
				if(in == 3) begin
					state<=7778;
					out<=199;
				end
				if(in == 4) begin
					state<=3889;
					out<=200;
				end
			end
			5877: begin
				if(in == 0) begin
					state<=4798;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=900;
					out<=203;
				end
				if(in == 3) begin
					state<=6165;
					out<=204;
				end
				if(in == 4) begin
					state<=2276;
					out<=205;
				end
			end
			5878: begin
				if(in == 0) begin
					state<=4799;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=901;
					out<=208;
				end
				if(in == 3) begin
					state<=6166;
					out<=209;
				end
				if(in == 4) begin
					state<=2277;
					out<=210;
				end
			end
			5879: begin
				if(in == 0) begin
					state<=4800;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=902;
					out<=213;
				end
				if(in == 3) begin
					state<=6167;
					out<=214;
				end
				if(in == 4) begin
					state<=2278;
					out<=215;
				end
			end
			5880: begin
				if(in == 0) begin
					state<=4801;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=903;
					out<=218;
				end
				if(in == 3) begin
					state<=6168;
					out<=219;
				end
				if(in == 4) begin
					state<=2279;
					out<=220;
				end
			end
			5881: begin
				if(in == 0) begin
					state<=4802;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=904;
					out<=223;
				end
				if(in == 3) begin
					state<=6169;
					out<=224;
				end
				if(in == 4) begin
					state<=2280;
					out<=225;
				end
			end
			5882: begin
				if(in == 0) begin
					state<=4803;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=905;
					out<=228;
				end
				if(in == 3) begin
					state<=6170;
					out<=229;
				end
				if(in == 4) begin
					state<=2281;
					out<=230;
				end
			end
			5883: begin
				if(in == 0) begin
					state<=4804;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=906;
					out<=233;
				end
				if(in == 3) begin
					state<=6171;
					out<=234;
				end
				if(in == 4) begin
					state<=2282;
					out<=235;
				end
			end
			5884: begin
				if(in == 0) begin
					state<=4805;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=907;
					out<=238;
				end
				if(in == 3) begin
					state<=6172;
					out<=239;
				end
				if(in == 4) begin
					state<=2283;
					out<=240;
				end
			end
			5885: begin
				if(in == 0) begin
					state<=4806;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=908;
					out<=243;
				end
				if(in == 3) begin
					state<=6173;
					out<=244;
				end
				if(in == 4) begin
					state<=2284;
					out<=245;
				end
			end
			5886: begin
				if(in == 0) begin
					state<=5887;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=1998;
					out<=248;
				end
				if(in == 3) begin
					state<=6164;
					out<=249;
				end
				if(in == 4) begin
					state<=2275;
					out<=250;
				end
			end
			5887: begin
				if(in == 0) begin
					state<=4808;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=910;
					out<=253;
				end
				if(in == 3) begin
					state<=6175;
					out<=254;
				end
				if(in == 4) begin
					state<=2286;
					out<=255;
				end
			end
			5888: begin
				if(in == 0) begin
					state<=5899;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=2010;
					out<=2;
				end
				if(in == 3) begin
					state<=3910;
					out<=3;
				end
				if(in == 4) begin
					state<=12;
					out<=4;
				end
			end
			5889: begin
				if(in == 0) begin
					state<=5900;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=2011;
					out<=7;
				end
				if(in == 3) begin
					state<=3911;
					out<=8;
				end
				if(in == 4) begin
					state<=13;
					out<=9;
				end
			end
			5890: begin
				if(in == 0) begin
					state<=5901;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=2012;
					out<=12;
				end
				if(in == 3) begin
					state<=3912;
					out<=13;
				end
				if(in == 4) begin
					state<=14;
					out<=14;
				end
			end
			5891: begin
				if(in == 0) begin
					state<=5902;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=2013;
					out<=17;
				end
				if(in == 3) begin
					state<=3913;
					out<=18;
				end
				if(in == 4) begin
					state<=15;
					out<=19;
				end
			end
			5892: begin
				if(in == 0) begin
					state<=5903;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=2014;
					out<=22;
				end
				if(in == 3) begin
					state<=3914;
					out<=23;
				end
				if(in == 4) begin
					state<=16;
					out<=24;
				end
			end
			5893: begin
				if(in == 0) begin
					state<=5904;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=2015;
					out<=27;
				end
				if(in == 3) begin
					state<=3915;
					out<=28;
				end
				if(in == 4) begin
					state<=17;
					out<=29;
				end
			end
			5894: begin
				if(in == 0) begin
					state<=5905;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=2016;
					out<=32;
				end
				if(in == 3) begin
					state<=3916;
					out<=33;
				end
				if(in == 4) begin
					state<=18;
					out<=34;
				end
			end
			5895: begin
				if(in == 0) begin
					state<=5906;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=2017;
					out<=37;
				end
				if(in == 3) begin
					state<=3917;
					out<=38;
				end
				if(in == 4) begin
					state<=19;
					out<=39;
				end
			end
			5896: begin
				if(in == 0) begin
					state<=5907;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=2018;
					out<=42;
				end
				if(in == 3) begin
					state<=3918;
					out<=43;
				end
				if(in == 4) begin
					state<=20;
					out<=44;
				end
			end
			5897: begin
				if(in == 0) begin
					state<=5898;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=2009;
					out<=47;
				end
				if(in == 3) begin
					state<=3909;
					out<=48;
				end
				if(in == 4) begin
					state<=11;
					out<=49;
				end
			end
			5898: begin
				if(in == 0) begin
					state<=5909;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=2020;
					out<=52;
				end
				if(in == 3) begin
					state<=3920;
					out<=53;
				end
				if(in == 4) begin
					state<=22;
					out<=54;
				end
			end
			5899: begin
				if(in == 0) begin
					state<=5910;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=2021;
					out<=57;
				end
				if(in == 3) begin
					state<=3921;
					out<=58;
				end
				if(in == 4) begin
					state<=23;
					out<=59;
				end
			end
			5900: begin
				if(in == 0) begin
					state<=5911;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=2022;
					out<=62;
				end
				if(in == 3) begin
					state<=3922;
					out<=63;
				end
				if(in == 4) begin
					state<=24;
					out<=64;
				end
			end
			5901: begin
				if(in == 0) begin
					state<=5912;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=2023;
					out<=67;
				end
				if(in == 3) begin
					state<=3923;
					out<=68;
				end
				if(in == 4) begin
					state<=25;
					out<=69;
				end
			end
			5902: begin
				if(in == 0) begin
					state<=5913;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=2024;
					out<=72;
				end
				if(in == 3) begin
					state<=3924;
					out<=73;
				end
				if(in == 4) begin
					state<=26;
					out<=74;
				end
			end
			5903: begin
				if(in == 0) begin
					state<=5914;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=2025;
					out<=77;
				end
				if(in == 3) begin
					state<=3925;
					out<=78;
				end
				if(in == 4) begin
					state<=27;
					out<=79;
				end
			end
			5904: begin
				if(in == 0) begin
					state<=5915;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=2026;
					out<=82;
				end
				if(in == 3) begin
					state<=3926;
					out<=83;
				end
				if(in == 4) begin
					state<=28;
					out<=84;
				end
			end
			5905: begin
				if(in == 0) begin
					state<=5916;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=2027;
					out<=87;
				end
				if(in == 3) begin
					state<=3927;
					out<=88;
				end
				if(in == 4) begin
					state<=29;
					out<=89;
				end
			end
			5906: begin
				if(in == 0) begin
					state<=5917;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=2028;
					out<=92;
				end
				if(in == 3) begin
					state<=3928;
					out<=93;
				end
				if(in == 4) begin
					state<=30;
					out<=94;
				end
			end
			5907: begin
				if(in == 0) begin
					state<=5908;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=2019;
					out<=97;
				end
				if(in == 3) begin
					state<=3919;
					out<=98;
				end
				if(in == 4) begin
					state<=21;
					out<=99;
				end
			end
			5908: begin
				if(in == 0) begin
					state<=5919;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=2030;
					out<=102;
				end
				if(in == 3) begin
					state<=3930;
					out<=103;
				end
				if(in == 4) begin
					state<=32;
					out<=104;
				end
			end
			5909: begin
				if(in == 0) begin
					state<=5920;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=2031;
					out<=107;
				end
				if(in == 3) begin
					state<=3931;
					out<=108;
				end
				if(in == 4) begin
					state<=33;
					out<=109;
				end
			end
			5910: begin
				if(in == 0) begin
					state<=5921;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=2032;
					out<=112;
				end
				if(in == 3) begin
					state<=3932;
					out<=113;
				end
				if(in == 4) begin
					state<=34;
					out<=114;
				end
			end
			5911: begin
				if(in == 0) begin
					state<=5922;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=2033;
					out<=117;
				end
				if(in == 3) begin
					state<=3933;
					out<=118;
				end
				if(in == 4) begin
					state<=35;
					out<=119;
				end
			end
			5912: begin
				if(in == 0) begin
					state<=5923;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=2034;
					out<=122;
				end
				if(in == 3) begin
					state<=3934;
					out<=123;
				end
				if(in == 4) begin
					state<=36;
					out<=124;
				end
			end
			5913: begin
				if(in == 0) begin
					state<=5924;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=2035;
					out<=127;
				end
				if(in == 3) begin
					state<=3935;
					out<=128;
				end
				if(in == 4) begin
					state<=37;
					out<=129;
				end
			end
			5914: begin
				if(in == 0) begin
					state<=5925;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=2036;
					out<=132;
				end
				if(in == 3) begin
					state<=3936;
					out<=133;
				end
				if(in == 4) begin
					state<=38;
					out<=134;
				end
			end
			5915: begin
				if(in == 0) begin
					state<=5926;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=2037;
					out<=137;
				end
				if(in == 3) begin
					state<=3937;
					out<=138;
				end
				if(in == 4) begin
					state<=39;
					out<=139;
				end
			end
			5916: begin
				if(in == 0) begin
					state<=5927;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=2038;
					out<=142;
				end
				if(in == 3) begin
					state<=3938;
					out<=143;
				end
				if(in == 4) begin
					state<=40;
					out<=144;
				end
			end
			5917: begin
				if(in == 0) begin
					state<=5918;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=2029;
					out<=147;
				end
				if(in == 3) begin
					state<=3929;
					out<=148;
				end
				if(in == 4) begin
					state<=31;
					out<=149;
				end
			end
			5918: begin
				if(in == 0) begin
					state<=5929;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=2040;
					out<=152;
				end
				if(in == 3) begin
					state<=3940;
					out<=153;
				end
				if(in == 4) begin
					state<=42;
					out<=154;
				end
			end
			5919: begin
				if(in == 0) begin
					state<=5930;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=2041;
					out<=157;
				end
				if(in == 3) begin
					state<=3941;
					out<=158;
				end
				if(in == 4) begin
					state<=43;
					out<=159;
				end
			end
			5920: begin
				if(in == 0) begin
					state<=5931;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=2042;
					out<=162;
				end
				if(in == 3) begin
					state<=3942;
					out<=163;
				end
				if(in == 4) begin
					state<=44;
					out<=164;
				end
			end
			5921: begin
				if(in == 0) begin
					state<=5932;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=2043;
					out<=167;
				end
				if(in == 3) begin
					state<=3943;
					out<=168;
				end
				if(in == 4) begin
					state<=45;
					out<=169;
				end
			end
			5922: begin
				if(in == 0) begin
					state<=5933;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=2044;
					out<=172;
				end
				if(in == 3) begin
					state<=3944;
					out<=173;
				end
				if(in == 4) begin
					state<=46;
					out<=174;
				end
			end
			5923: begin
				if(in == 0) begin
					state<=5934;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=2045;
					out<=177;
				end
				if(in == 3) begin
					state<=3945;
					out<=178;
				end
				if(in == 4) begin
					state<=47;
					out<=179;
				end
			end
			5924: begin
				if(in == 0) begin
					state<=5935;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=2046;
					out<=182;
				end
				if(in == 3) begin
					state<=3946;
					out<=183;
				end
				if(in == 4) begin
					state<=48;
					out<=184;
				end
			end
			5925: begin
				if(in == 0) begin
					state<=5936;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=2047;
					out<=187;
				end
				if(in == 3) begin
					state<=3947;
					out<=188;
				end
				if(in == 4) begin
					state<=49;
					out<=189;
				end
			end
			5926: begin
				if(in == 0) begin
					state<=5937;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=2048;
					out<=192;
				end
				if(in == 3) begin
					state<=3948;
					out<=193;
				end
				if(in == 4) begin
					state<=50;
					out<=194;
				end
			end
			5927: begin
				if(in == 0) begin
					state<=5928;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=2039;
					out<=197;
				end
				if(in == 3) begin
					state<=3939;
					out<=198;
				end
				if(in == 4) begin
					state<=41;
					out<=199;
				end
			end
			5928: begin
				if(in == 0) begin
					state<=7151;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=3262;
					out<=202;
				end
				if(in == 3) begin
					state<=5219;
					out<=203;
				end
				if(in == 4) begin
					state<=1330;
					out<=204;
				end
			end
			5929: begin
				if(in == 0) begin
					state<=7152;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=3263;
					out<=207;
				end
				if(in == 3) begin
					state<=5220;
					out<=208;
				end
				if(in == 4) begin
					state<=1331;
					out<=209;
				end
			end
			5930: begin
				if(in == 0) begin
					state<=7153;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=3264;
					out<=212;
				end
				if(in == 3) begin
					state<=5221;
					out<=213;
				end
				if(in == 4) begin
					state<=1332;
					out<=214;
				end
			end
			5931: begin
				if(in == 0) begin
					state<=7154;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=3265;
					out<=217;
				end
				if(in == 3) begin
					state<=5222;
					out<=218;
				end
				if(in == 4) begin
					state<=1333;
					out<=219;
				end
			end
			5932: begin
				if(in == 0) begin
					state<=7155;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=3266;
					out<=222;
				end
				if(in == 3) begin
					state<=5223;
					out<=223;
				end
				if(in == 4) begin
					state<=1334;
					out<=224;
				end
			end
			5933: begin
				if(in == 0) begin
					state<=7156;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=3267;
					out<=227;
				end
				if(in == 3) begin
					state<=5224;
					out<=228;
				end
				if(in == 4) begin
					state<=1335;
					out<=229;
				end
			end
			5934: begin
				if(in == 0) begin
					state<=7157;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=3268;
					out<=232;
				end
				if(in == 3) begin
					state<=5225;
					out<=233;
				end
				if(in == 4) begin
					state<=1336;
					out<=234;
				end
			end
			5935: begin
				if(in == 0) begin
					state<=7158;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=3269;
					out<=237;
				end
				if(in == 3) begin
					state<=5226;
					out<=238;
				end
				if(in == 4) begin
					state<=1337;
					out<=239;
				end
			end
			5936: begin
				if(in == 0) begin
					state<=7159;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=3270;
					out<=242;
				end
				if(in == 3) begin
					state<=5227;
					out<=243;
				end
				if(in == 4) begin
					state<=1338;
					out<=244;
				end
			end
			5937: begin
				if(in == 0) begin
					state<=7150;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=3261;
					out<=247;
				end
				if(in == 3) begin
					state<=5218;
					out<=248;
				end
				if(in == 4) begin
					state<=1329;
					out<=249;
				end
			end
			5938: begin
				if(in == 0) begin
					state<=5949;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=2060;
					out<=252;
				end
				if(in == 3) begin
					state<=3960;
					out<=253;
				end
				if(in == 4) begin
					state<=62;
					out<=254;
				end
			end
			5939: begin
				if(in == 0) begin
					state<=5950;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=2061;
					out<=1;
				end
				if(in == 3) begin
					state<=3961;
					out<=2;
				end
				if(in == 4) begin
					state<=63;
					out<=3;
				end
			end
			5940: begin
				if(in == 0) begin
					state<=5951;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=2062;
					out<=6;
				end
				if(in == 3) begin
					state<=3962;
					out<=7;
				end
				if(in == 4) begin
					state<=64;
					out<=8;
				end
			end
			5941: begin
				if(in == 0) begin
					state<=5952;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=2063;
					out<=11;
				end
				if(in == 3) begin
					state<=3963;
					out<=12;
				end
				if(in == 4) begin
					state<=65;
					out<=13;
				end
			end
			5942: begin
				if(in == 0) begin
					state<=5953;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=2064;
					out<=16;
				end
				if(in == 3) begin
					state<=3964;
					out<=17;
				end
				if(in == 4) begin
					state<=66;
					out<=18;
				end
			end
			5943: begin
				if(in == 0) begin
					state<=5954;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=2065;
					out<=21;
				end
				if(in == 3) begin
					state<=3965;
					out<=22;
				end
				if(in == 4) begin
					state<=67;
					out<=23;
				end
			end
			5944: begin
				if(in == 0) begin
					state<=5955;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=2066;
					out<=26;
				end
				if(in == 3) begin
					state<=3966;
					out<=27;
				end
				if(in == 4) begin
					state<=68;
					out<=28;
				end
			end
			5945: begin
				if(in == 0) begin
					state<=5956;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=2067;
					out<=31;
				end
				if(in == 3) begin
					state<=3967;
					out<=32;
				end
				if(in == 4) begin
					state<=69;
					out<=33;
				end
			end
			5946: begin
				if(in == 0) begin
					state<=5947;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=2058;
					out<=36;
				end
				if(in == 3) begin
					state<=3958;
					out<=37;
				end
				if(in == 4) begin
					state<=60;
					out<=38;
				end
			end
			5947: begin
				if(in == 0) begin
					state<=5958;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=2069;
					out<=41;
				end
				if(in == 3) begin
					state<=3969;
					out<=42;
				end
				if(in == 4) begin
					state<=71;
					out<=43;
				end
			end
			5948: begin
				if(in == 0) begin
					state<=5959;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=2070;
					out<=46;
				end
				if(in == 3) begin
					state<=3970;
					out<=47;
				end
				if(in == 4) begin
					state<=72;
					out<=48;
				end
			end
			5949: begin
				if(in == 0) begin
					state<=5960;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=2071;
					out<=51;
				end
				if(in == 3) begin
					state<=3971;
					out<=52;
				end
				if(in == 4) begin
					state<=73;
					out<=53;
				end
			end
			5950: begin
				if(in == 0) begin
					state<=5961;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=2072;
					out<=56;
				end
				if(in == 3) begin
					state<=3972;
					out<=57;
				end
				if(in == 4) begin
					state<=74;
					out<=58;
				end
			end
			5951: begin
				if(in == 0) begin
					state<=5962;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=2073;
					out<=61;
				end
				if(in == 3) begin
					state<=3973;
					out<=62;
				end
				if(in == 4) begin
					state<=75;
					out<=63;
				end
			end
			5952: begin
				if(in == 0) begin
					state<=5963;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=2074;
					out<=66;
				end
				if(in == 3) begin
					state<=3974;
					out<=67;
				end
				if(in == 4) begin
					state<=76;
					out<=68;
				end
			end
			5953: begin
				if(in == 0) begin
					state<=5964;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=2075;
					out<=71;
				end
				if(in == 3) begin
					state<=3975;
					out<=72;
				end
				if(in == 4) begin
					state<=77;
					out<=73;
				end
			end
			5954: begin
				if(in == 0) begin
					state<=5965;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=2076;
					out<=76;
				end
				if(in == 3) begin
					state<=3976;
					out<=77;
				end
				if(in == 4) begin
					state<=78;
					out<=78;
				end
			end
			5955: begin
				if(in == 0) begin
					state<=5966;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=2077;
					out<=81;
				end
				if(in == 3) begin
					state<=3977;
					out<=82;
				end
				if(in == 4) begin
					state<=79;
					out<=83;
				end
			end
			5956: begin
				if(in == 0) begin
					state<=5957;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=2068;
					out<=86;
				end
				if(in == 3) begin
					state<=3968;
					out<=87;
				end
				if(in == 4) begin
					state<=70;
					out<=88;
				end
			end
			5957: begin
				if(in == 0) begin
					state<=5968;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=2079;
					out<=91;
				end
				if(in == 3) begin
					state<=3979;
					out<=92;
				end
				if(in == 4) begin
					state<=81;
					out<=93;
				end
			end
			5958: begin
				if(in == 0) begin
					state<=5969;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=2080;
					out<=96;
				end
				if(in == 3) begin
					state<=3980;
					out<=97;
				end
				if(in == 4) begin
					state<=82;
					out<=98;
				end
			end
			5959: begin
				if(in == 0) begin
					state<=5970;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=2081;
					out<=101;
				end
				if(in == 3) begin
					state<=3981;
					out<=102;
				end
				if(in == 4) begin
					state<=83;
					out<=103;
				end
			end
			5960: begin
				if(in == 0) begin
					state<=5971;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=2082;
					out<=106;
				end
				if(in == 3) begin
					state<=3982;
					out<=107;
				end
				if(in == 4) begin
					state<=84;
					out<=108;
				end
			end
			5961: begin
				if(in == 0) begin
					state<=5972;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=2083;
					out<=111;
				end
				if(in == 3) begin
					state<=3983;
					out<=112;
				end
				if(in == 4) begin
					state<=85;
					out<=113;
				end
			end
			5962: begin
				if(in == 0) begin
					state<=5973;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=2084;
					out<=116;
				end
				if(in == 3) begin
					state<=3984;
					out<=117;
				end
				if(in == 4) begin
					state<=86;
					out<=118;
				end
			end
			5963: begin
				if(in == 0) begin
					state<=5974;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=2085;
					out<=121;
				end
				if(in == 3) begin
					state<=3985;
					out<=122;
				end
				if(in == 4) begin
					state<=87;
					out<=123;
				end
			end
			5964: begin
				if(in == 0) begin
					state<=5975;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=2086;
					out<=126;
				end
				if(in == 3) begin
					state<=3986;
					out<=127;
				end
				if(in == 4) begin
					state<=88;
					out<=128;
				end
			end
			5965: begin
				if(in == 0) begin
					state<=5976;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=2087;
					out<=131;
				end
				if(in == 3) begin
					state<=3987;
					out<=132;
				end
				if(in == 4) begin
					state<=89;
					out<=133;
				end
			end
			5966: begin
				if(in == 0) begin
					state<=5967;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=2078;
					out<=136;
				end
				if(in == 3) begin
					state<=3978;
					out<=137;
				end
				if(in == 4) begin
					state<=80;
					out<=138;
				end
			end
			5967: begin
				if(in == 0) begin
					state<=5978;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=2089;
					out<=141;
				end
				if(in == 3) begin
					state<=3989;
					out<=142;
				end
				if(in == 4) begin
					state<=91;
					out<=143;
				end
			end
			5968: begin
				if(in == 0) begin
					state<=5979;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=2090;
					out<=146;
				end
				if(in == 3) begin
					state<=3990;
					out<=147;
				end
				if(in == 4) begin
					state<=92;
					out<=148;
				end
			end
			5969: begin
				if(in == 0) begin
					state<=5980;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=2091;
					out<=151;
				end
				if(in == 3) begin
					state<=3991;
					out<=152;
				end
				if(in == 4) begin
					state<=93;
					out<=153;
				end
			end
			5970: begin
				if(in == 0) begin
					state<=5981;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=2092;
					out<=156;
				end
				if(in == 3) begin
					state<=3992;
					out<=157;
				end
				if(in == 4) begin
					state<=94;
					out<=158;
				end
			end
			5971: begin
				if(in == 0) begin
					state<=5982;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=2093;
					out<=161;
				end
				if(in == 3) begin
					state<=3993;
					out<=162;
				end
				if(in == 4) begin
					state<=95;
					out<=163;
				end
			end
			5972: begin
				if(in == 0) begin
					state<=5983;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=2094;
					out<=166;
				end
				if(in == 3) begin
					state<=3994;
					out<=167;
				end
				if(in == 4) begin
					state<=96;
					out<=168;
				end
			end
			5973: begin
				if(in == 0) begin
					state<=5984;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=2095;
					out<=171;
				end
				if(in == 3) begin
					state<=3995;
					out<=172;
				end
				if(in == 4) begin
					state<=97;
					out<=173;
				end
			end
			5974: begin
				if(in == 0) begin
					state<=5985;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=2096;
					out<=176;
				end
				if(in == 3) begin
					state<=3996;
					out<=177;
				end
				if(in == 4) begin
					state<=98;
					out<=178;
				end
			end
			5975: begin
				if(in == 0) begin
					state<=5986;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=2097;
					out<=181;
				end
				if(in == 3) begin
					state<=3997;
					out<=182;
				end
				if(in == 4) begin
					state<=99;
					out<=183;
				end
			end
			5976: begin
				if(in == 0) begin
					state<=5977;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=2088;
					out<=186;
				end
				if(in == 3) begin
					state<=3988;
					out<=187;
				end
				if(in == 4) begin
					state<=90;
					out<=188;
				end
			end
			5977: begin
				if(in == 0) begin
					state<=5988;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=2099;
					out<=191;
				end
				if(in == 3) begin
					state<=3999;
					out<=192;
				end
				if(in == 4) begin
					state<=101;
					out<=193;
				end
			end
			5978: begin
				if(in == 0) begin
					state<=5989;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=2100;
					out<=196;
				end
				if(in == 3) begin
					state<=4000;
					out<=197;
				end
				if(in == 4) begin
					state<=102;
					out<=198;
				end
			end
			5979: begin
				if(in == 0) begin
					state<=5990;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=2101;
					out<=201;
				end
				if(in == 3) begin
					state<=4001;
					out<=202;
				end
				if(in == 4) begin
					state<=103;
					out<=203;
				end
			end
			5980: begin
				if(in == 0) begin
					state<=5991;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=2102;
					out<=206;
				end
				if(in == 3) begin
					state<=4002;
					out<=207;
				end
				if(in == 4) begin
					state<=104;
					out<=208;
				end
			end
			5981: begin
				if(in == 0) begin
					state<=5992;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=2103;
					out<=211;
				end
				if(in == 3) begin
					state<=4003;
					out<=212;
				end
				if(in == 4) begin
					state<=105;
					out<=213;
				end
			end
			5982: begin
				if(in == 0) begin
					state<=5993;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=2104;
					out<=216;
				end
				if(in == 3) begin
					state<=4004;
					out<=217;
				end
				if(in == 4) begin
					state<=106;
					out<=218;
				end
			end
			5983: begin
				if(in == 0) begin
					state<=5994;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=2105;
					out<=221;
				end
				if(in == 3) begin
					state<=4005;
					out<=222;
				end
				if(in == 4) begin
					state<=107;
					out<=223;
				end
			end
			5984: begin
				if(in == 0) begin
					state<=5995;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=2106;
					out<=226;
				end
				if(in == 3) begin
					state<=4006;
					out<=227;
				end
				if(in == 4) begin
					state<=108;
					out<=228;
				end
			end
			5985: begin
				if(in == 0) begin
					state<=5996;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=2107;
					out<=231;
				end
				if(in == 3) begin
					state<=4007;
					out<=232;
				end
				if(in == 4) begin
					state<=109;
					out<=233;
				end
			end
			5986: begin
				if(in == 0) begin
					state<=5987;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=2098;
					out<=236;
				end
				if(in == 3) begin
					state<=3998;
					out<=237;
				end
				if(in == 4) begin
					state<=100;
					out<=238;
				end
			end
			5987: begin
				if(in == 0) begin
					state<=5998;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=2109;
					out<=241;
				end
				if(in == 3) begin
					state<=4009;
					out<=242;
				end
				if(in == 4) begin
					state<=111;
					out<=243;
				end
			end
			5988: begin
				if(in == 0) begin
					state<=5999;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=2110;
					out<=246;
				end
				if(in == 3) begin
					state<=4010;
					out<=247;
				end
				if(in == 4) begin
					state<=112;
					out<=248;
				end
			end
			5989: begin
				if(in == 0) begin
					state<=6000;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=2111;
					out<=251;
				end
				if(in == 3) begin
					state<=4011;
					out<=252;
				end
				if(in == 4) begin
					state<=113;
					out<=253;
				end
			end
			5990: begin
				if(in == 0) begin
					state<=6001;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=2112;
					out<=0;
				end
				if(in == 3) begin
					state<=4012;
					out<=1;
				end
				if(in == 4) begin
					state<=114;
					out<=2;
				end
			end
			5991: begin
				if(in == 0) begin
					state<=6002;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=2113;
					out<=5;
				end
				if(in == 3) begin
					state<=4013;
					out<=6;
				end
				if(in == 4) begin
					state<=115;
					out<=7;
				end
			end
			5992: begin
				if(in == 0) begin
					state<=6003;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=2114;
					out<=10;
				end
				if(in == 3) begin
					state<=4014;
					out<=11;
				end
				if(in == 4) begin
					state<=116;
					out<=12;
				end
			end
			5993: begin
				if(in == 0) begin
					state<=6004;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=2115;
					out<=15;
				end
				if(in == 3) begin
					state<=4015;
					out<=16;
				end
				if(in == 4) begin
					state<=117;
					out<=17;
				end
			end
			5994: begin
				if(in == 0) begin
					state<=6005;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=2116;
					out<=20;
				end
				if(in == 3) begin
					state<=4016;
					out<=21;
				end
				if(in == 4) begin
					state<=118;
					out<=22;
				end
			end
			5995: begin
				if(in == 0) begin
					state<=6006;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=2117;
					out<=25;
				end
				if(in == 3) begin
					state<=4017;
					out<=26;
				end
				if(in == 4) begin
					state<=119;
					out<=27;
				end
			end
			5996: begin
				if(in == 0) begin
					state<=5997;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=2108;
					out<=30;
				end
				if(in == 3) begin
					state<=4008;
					out<=31;
				end
				if(in == 4) begin
					state<=110;
					out<=32;
				end
			end
			5997: begin
				if(in == 0) begin
					state<=7182;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=3293;
					out<=35;
				end
				if(in == 3) begin
					state<=5250;
					out<=36;
				end
				if(in == 4) begin
					state<=1361;
					out<=37;
				end
			end
			5998: begin
				if(in == 0) begin
					state<=7183;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=3294;
					out<=40;
				end
				if(in == 3) begin
					state<=5251;
					out<=41;
				end
				if(in == 4) begin
					state<=1362;
					out<=42;
				end
			end
			5999: begin
				if(in == 0) begin
					state<=7184;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=3295;
					out<=45;
				end
				if(in == 3) begin
					state<=5252;
					out<=46;
				end
				if(in == 4) begin
					state<=1363;
					out<=47;
				end
			end
			6000: begin
				if(in == 0) begin
					state<=7185;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=3296;
					out<=50;
				end
				if(in == 3) begin
					state<=5253;
					out<=51;
				end
				if(in == 4) begin
					state<=1364;
					out<=52;
				end
			end
			6001: begin
				if(in == 0) begin
					state<=7186;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=3297;
					out<=55;
				end
				if(in == 3) begin
					state<=5254;
					out<=56;
				end
				if(in == 4) begin
					state<=1365;
					out<=57;
				end
			end
			6002: begin
				if(in == 0) begin
					state<=7187;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=3298;
					out<=60;
				end
				if(in == 3) begin
					state<=5255;
					out<=61;
				end
				if(in == 4) begin
					state<=1366;
					out<=62;
				end
			end
			6003: begin
				if(in == 0) begin
					state<=7188;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=3299;
					out<=65;
				end
				if(in == 3) begin
					state<=5256;
					out<=66;
				end
				if(in == 4) begin
					state<=1367;
					out<=67;
				end
			end
			6004: begin
				if(in == 0) begin
					state<=7189;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=3300;
					out<=70;
				end
				if(in == 3) begin
					state<=5257;
					out<=71;
				end
				if(in == 4) begin
					state<=1368;
					out<=72;
				end
			end
			6005: begin
				if(in == 0) begin
					state<=7190;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=3301;
					out<=75;
				end
				if(in == 3) begin
					state<=5258;
					out<=76;
				end
				if(in == 4) begin
					state<=1369;
					out<=77;
				end
			end
			6006: begin
				if(in == 0) begin
					state<=7181;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=3292;
					out<=80;
				end
				if(in == 3) begin
					state<=5249;
					out<=81;
				end
				if(in == 4) begin
					state<=1360;
					out<=82;
				end
			end
			6007: begin
				if(in == 0) begin
					state<=6018;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=2129;
					out<=85;
				end
				if(in == 3) begin
					state<=4029;
					out<=86;
				end
				if(in == 4) begin
					state<=131;
					out<=87;
				end
			end
			6008: begin
				if(in == 0) begin
					state<=6019;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=2130;
					out<=90;
				end
				if(in == 3) begin
					state<=4030;
					out<=91;
				end
				if(in == 4) begin
					state<=132;
					out<=92;
				end
			end
			6009: begin
				if(in == 0) begin
					state<=6020;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=2131;
					out<=95;
				end
				if(in == 3) begin
					state<=4031;
					out<=96;
				end
				if(in == 4) begin
					state<=133;
					out<=97;
				end
			end
			6010: begin
				if(in == 0) begin
					state<=6021;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=2132;
					out<=100;
				end
				if(in == 3) begin
					state<=4032;
					out<=101;
				end
				if(in == 4) begin
					state<=134;
					out<=102;
				end
			end
			6011: begin
				if(in == 0) begin
					state<=6022;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=2133;
					out<=105;
				end
				if(in == 3) begin
					state<=4033;
					out<=106;
				end
				if(in == 4) begin
					state<=135;
					out<=107;
				end
			end
			6012: begin
				if(in == 0) begin
					state<=6023;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=2134;
					out<=110;
				end
				if(in == 3) begin
					state<=4034;
					out<=111;
				end
				if(in == 4) begin
					state<=136;
					out<=112;
				end
			end
			6013: begin
				if(in == 0) begin
					state<=6024;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=2135;
					out<=115;
				end
				if(in == 3) begin
					state<=4035;
					out<=116;
				end
				if(in == 4) begin
					state<=137;
					out<=117;
				end
			end
			6014: begin
				if(in == 0) begin
					state<=6025;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=2136;
					out<=120;
				end
				if(in == 3) begin
					state<=4036;
					out<=121;
				end
				if(in == 4) begin
					state<=138;
					out<=122;
				end
			end
			6015: begin
				if(in == 0) begin
					state<=6016;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=2127;
					out<=125;
				end
				if(in == 3) begin
					state<=4027;
					out<=126;
				end
				if(in == 4) begin
					state<=129;
					out<=127;
				end
			end
			6016: begin
				if(in == 0) begin
					state<=6027;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=2138;
					out<=130;
				end
				if(in == 3) begin
					state<=4038;
					out<=131;
				end
				if(in == 4) begin
					state<=140;
					out<=132;
				end
			end
			6017: begin
				if(in == 0) begin
					state<=6028;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=2139;
					out<=135;
				end
				if(in == 3) begin
					state<=4039;
					out<=136;
				end
				if(in == 4) begin
					state<=141;
					out<=137;
				end
			end
			6018: begin
				if(in == 0) begin
					state<=6029;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=2140;
					out<=140;
				end
				if(in == 3) begin
					state<=4040;
					out<=141;
				end
				if(in == 4) begin
					state<=142;
					out<=142;
				end
			end
			6019: begin
				if(in == 0) begin
					state<=6030;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=2141;
					out<=145;
				end
				if(in == 3) begin
					state<=4041;
					out<=146;
				end
				if(in == 4) begin
					state<=143;
					out<=147;
				end
			end
			6020: begin
				if(in == 0) begin
					state<=6031;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=2142;
					out<=150;
				end
				if(in == 3) begin
					state<=4042;
					out<=151;
				end
				if(in == 4) begin
					state<=144;
					out<=152;
				end
			end
			6021: begin
				if(in == 0) begin
					state<=6032;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=2143;
					out<=155;
				end
				if(in == 3) begin
					state<=4043;
					out<=156;
				end
				if(in == 4) begin
					state<=145;
					out<=157;
				end
			end
			6022: begin
				if(in == 0) begin
					state<=6033;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=2144;
					out<=160;
				end
				if(in == 3) begin
					state<=4044;
					out<=161;
				end
				if(in == 4) begin
					state<=146;
					out<=162;
				end
			end
			6023: begin
				if(in == 0) begin
					state<=6034;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=2145;
					out<=165;
				end
				if(in == 3) begin
					state<=4045;
					out<=166;
				end
				if(in == 4) begin
					state<=147;
					out<=167;
				end
			end
			6024: begin
				if(in == 0) begin
					state<=6035;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=2146;
					out<=170;
				end
				if(in == 3) begin
					state<=4046;
					out<=171;
				end
				if(in == 4) begin
					state<=148;
					out<=172;
				end
			end
			6025: begin
				if(in == 0) begin
					state<=6026;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=2137;
					out<=175;
				end
				if(in == 3) begin
					state<=4037;
					out<=176;
				end
				if(in == 4) begin
					state<=139;
					out<=177;
				end
			end
			6026: begin
				if(in == 0) begin
					state<=6037;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=2148;
					out<=180;
				end
				if(in == 3) begin
					state<=4048;
					out<=181;
				end
				if(in == 4) begin
					state<=150;
					out<=182;
				end
			end
			6027: begin
				if(in == 0) begin
					state<=6038;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=2149;
					out<=185;
				end
				if(in == 3) begin
					state<=4049;
					out<=186;
				end
				if(in == 4) begin
					state<=151;
					out<=187;
				end
			end
			6028: begin
				if(in == 0) begin
					state<=6039;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=2150;
					out<=190;
				end
				if(in == 3) begin
					state<=4050;
					out<=191;
				end
				if(in == 4) begin
					state<=152;
					out<=192;
				end
			end
			6029: begin
				if(in == 0) begin
					state<=6040;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=2151;
					out<=195;
				end
				if(in == 3) begin
					state<=4051;
					out<=196;
				end
				if(in == 4) begin
					state<=153;
					out<=197;
				end
			end
			6030: begin
				if(in == 0) begin
					state<=6041;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=2152;
					out<=200;
				end
				if(in == 3) begin
					state<=4052;
					out<=201;
				end
				if(in == 4) begin
					state<=154;
					out<=202;
				end
			end
			6031: begin
				if(in == 0) begin
					state<=6042;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=2153;
					out<=205;
				end
				if(in == 3) begin
					state<=4053;
					out<=206;
				end
				if(in == 4) begin
					state<=155;
					out<=207;
				end
			end
			6032: begin
				if(in == 0) begin
					state<=6043;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=2154;
					out<=210;
				end
				if(in == 3) begin
					state<=4054;
					out<=211;
				end
				if(in == 4) begin
					state<=156;
					out<=212;
				end
			end
			6033: begin
				if(in == 0) begin
					state<=6044;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=2155;
					out<=215;
				end
				if(in == 3) begin
					state<=4055;
					out<=216;
				end
				if(in == 4) begin
					state<=157;
					out<=217;
				end
			end
			6034: begin
				if(in == 0) begin
					state<=6045;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=2156;
					out<=220;
				end
				if(in == 3) begin
					state<=4056;
					out<=221;
				end
				if(in == 4) begin
					state<=158;
					out<=222;
				end
			end
			6035: begin
				if(in == 0) begin
					state<=6036;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=2147;
					out<=225;
				end
				if(in == 3) begin
					state<=4047;
					out<=226;
				end
				if(in == 4) begin
					state<=149;
					out<=227;
				end
			end
			6036: begin
				if(in == 0) begin
					state<=6047;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=2158;
					out<=230;
				end
				if(in == 3) begin
					state<=4058;
					out<=231;
				end
				if(in == 4) begin
					state<=160;
					out<=232;
				end
			end
			6037: begin
				if(in == 0) begin
					state<=6048;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=2159;
					out<=235;
				end
				if(in == 3) begin
					state<=4059;
					out<=236;
				end
				if(in == 4) begin
					state<=161;
					out<=237;
				end
			end
			6038: begin
				if(in == 0) begin
					state<=6049;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=2160;
					out<=240;
				end
				if(in == 3) begin
					state<=4060;
					out<=241;
				end
				if(in == 4) begin
					state<=162;
					out<=242;
				end
			end
			6039: begin
				if(in == 0) begin
					state<=6050;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=2161;
					out<=245;
				end
				if(in == 3) begin
					state<=4061;
					out<=246;
				end
				if(in == 4) begin
					state<=163;
					out<=247;
				end
			end
			6040: begin
				if(in == 0) begin
					state<=6051;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=2162;
					out<=250;
				end
				if(in == 3) begin
					state<=4062;
					out<=251;
				end
				if(in == 4) begin
					state<=164;
					out<=252;
				end
			end
			6041: begin
				if(in == 0) begin
					state<=6052;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=2163;
					out<=255;
				end
				if(in == 3) begin
					state<=4063;
					out<=0;
				end
				if(in == 4) begin
					state<=165;
					out<=1;
				end
			end
			6042: begin
				if(in == 0) begin
					state<=6053;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=2164;
					out<=4;
				end
				if(in == 3) begin
					state<=4064;
					out<=5;
				end
				if(in == 4) begin
					state<=166;
					out<=6;
				end
			end
			6043: begin
				if(in == 0) begin
					state<=6054;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=2165;
					out<=9;
				end
				if(in == 3) begin
					state<=4065;
					out<=10;
				end
				if(in == 4) begin
					state<=167;
					out<=11;
				end
			end
			6044: begin
				if(in == 0) begin
					state<=6055;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=2166;
					out<=14;
				end
				if(in == 3) begin
					state<=4066;
					out<=15;
				end
				if(in == 4) begin
					state<=168;
					out<=16;
				end
			end
			6045: begin
				if(in == 0) begin
					state<=6046;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=2157;
					out<=19;
				end
				if(in == 3) begin
					state<=4057;
					out<=20;
				end
				if(in == 4) begin
					state<=159;
					out<=21;
				end
			end
			6046: begin
				if(in == 0) begin
					state<=6057;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=2168;
					out<=24;
				end
				if(in == 3) begin
					state<=4068;
					out<=25;
				end
				if(in == 4) begin
					state<=170;
					out<=26;
				end
			end
			6047: begin
				if(in == 0) begin
					state<=6058;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=2169;
					out<=29;
				end
				if(in == 3) begin
					state<=4069;
					out<=30;
				end
				if(in == 4) begin
					state<=171;
					out<=31;
				end
			end
			6048: begin
				if(in == 0) begin
					state<=6059;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=2170;
					out<=34;
				end
				if(in == 3) begin
					state<=4070;
					out<=35;
				end
				if(in == 4) begin
					state<=172;
					out<=36;
				end
			end
			6049: begin
				if(in == 0) begin
					state<=6060;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=2171;
					out<=39;
				end
				if(in == 3) begin
					state<=4071;
					out<=40;
				end
				if(in == 4) begin
					state<=173;
					out<=41;
				end
			end
			6050: begin
				if(in == 0) begin
					state<=6061;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=2172;
					out<=44;
				end
				if(in == 3) begin
					state<=4072;
					out<=45;
				end
				if(in == 4) begin
					state<=174;
					out<=46;
				end
			end
			6051: begin
				if(in == 0) begin
					state<=6062;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=2173;
					out<=49;
				end
				if(in == 3) begin
					state<=4073;
					out<=50;
				end
				if(in == 4) begin
					state<=175;
					out<=51;
				end
			end
			6052: begin
				if(in == 0) begin
					state<=6063;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=2174;
					out<=54;
				end
				if(in == 3) begin
					state<=4074;
					out<=55;
				end
				if(in == 4) begin
					state<=176;
					out<=56;
				end
			end
			6053: begin
				if(in == 0) begin
					state<=6064;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=2175;
					out<=59;
				end
				if(in == 3) begin
					state<=4075;
					out<=60;
				end
				if(in == 4) begin
					state<=177;
					out<=61;
				end
			end
			6054: begin
				if(in == 0) begin
					state<=6065;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=2176;
					out<=64;
				end
				if(in == 3) begin
					state<=4076;
					out<=65;
				end
				if(in == 4) begin
					state<=178;
					out<=66;
				end
			end
			6055: begin
				if(in == 0) begin
					state<=6056;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=2167;
					out<=69;
				end
				if(in == 3) begin
					state<=4067;
					out<=70;
				end
				if(in == 4) begin
					state<=169;
					out<=71;
				end
			end
			6056: begin
				if(in == 0) begin
					state<=6067;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=2178;
					out<=74;
				end
				if(in == 3) begin
					state<=4078;
					out<=75;
				end
				if(in == 4) begin
					state<=180;
					out<=76;
				end
			end
			6057: begin
				if(in == 0) begin
					state<=6068;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=2179;
					out<=79;
				end
				if(in == 3) begin
					state<=4079;
					out<=80;
				end
				if(in == 4) begin
					state<=181;
					out<=81;
				end
			end
			6058: begin
				if(in == 0) begin
					state<=6069;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=2180;
					out<=84;
				end
				if(in == 3) begin
					state<=4080;
					out<=85;
				end
				if(in == 4) begin
					state<=182;
					out<=86;
				end
			end
			6059: begin
				if(in == 0) begin
					state<=6070;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=2181;
					out<=89;
				end
				if(in == 3) begin
					state<=4081;
					out<=90;
				end
				if(in == 4) begin
					state<=183;
					out<=91;
				end
			end
			6060: begin
				if(in == 0) begin
					state<=6071;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=2182;
					out<=94;
				end
				if(in == 3) begin
					state<=4082;
					out<=95;
				end
				if(in == 4) begin
					state<=184;
					out<=96;
				end
			end
			6061: begin
				if(in == 0) begin
					state<=6072;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=2183;
					out<=99;
				end
				if(in == 3) begin
					state<=4083;
					out<=100;
				end
				if(in == 4) begin
					state<=185;
					out<=101;
				end
			end
			6062: begin
				if(in == 0) begin
					state<=6073;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=2184;
					out<=104;
				end
				if(in == 3) begin
					state<=4084;
					out<=105;
				end
				if(in == 4) begin
					state<=186;
					out<=106;
				end
			end
			6063: begin
				if(in == 0) begin
					state<=6074;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=2185;
					out<=109;
				end
				if(in == 3) begin
					state<=4085;
					out<=110;
				end
				if(in == 4) begin
					state<=187;
					out<=111;
				end
			end
			6064: begin
				if(in == 0) begin
					state<=6075;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=2186;
					out<=114;
				end
				if(in == 3) begin
					state<=4086;
					out<=115;
				end
				if(in == 4) begin
					state<=188;
					out<=116;
				end
			end
			6065: begin
				if(in == 0) begin
					state<=6066;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=2177;
					out<=119;
				end
				if(in == 3) begin
					state<=4077;
					out<=120;
				end
				if(in == 4) begin
					state<=179;
					out<=121;
				end
			end
			6066: begin
				if(in == 0) begin
					state<=7213;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=3324;
					out<=124;
				end
				if(in == 3) begin
					state<=5281;
					out<=125;
				end
				if(in == 4) begin
					state<=1392;
					out<=126;
				end
			end
			6067: begin
				if(in == 0) begin
					state<=7214;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=3325;
					out<=129;
				end
				if(in == 3) begin
					state<=5282;
					out<=130;
				end
				if(in == 4) begin
					state<=1393;
					out<=131;
				end
			end
			6068: begin
				if(in == 0) begin
					state<=7215;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=3326;
					out<=134;
				end
				if(in == 3) begin
					state<=5283;
					out<=135;
				end
				if(in == 4) begin
					state<=1394;
					out<=136;
				end
			end
			6069: begin
				if(in == 0) begin
					state<=7216;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=3327;
					out<=139;
				end
				if(in == 3) begin
					state<=5284;
					out<=140;
				end
				if(in == 4) begin
					state<=1395;
					out<=141;
				end
			end
			6070: begin
				if(in == 0) begin
					state<=7217;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=3328;
					out<=144;
				end
				if(in == 3) begin
					state<=5285;
					out<=145;
				end
				if(in == 4) begin
					state<=1396;
					out<=146;
				end
			end
			6071: begin
				if(in == 0) begin
					state<=7218;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=3329;
					out<=149;
				end
				if(in == 3) begin
					state<=5286;
					out<=150;
				end
				if(in == 4) begin
					state<=1397;
					out<=151;
				end
			end
			6072: begin
				if(in == 0) begin
					state<=7219;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=3330;
					out<=154;
				end
				if(in == 3) begin
					state<=5287;
					out<=155;
				end
				if(in == 4) begin
					state<=1398;
					out<=156;
				end
			end
			6073: begin
				if(in == 0) begin
					state<=7220;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=3331;
					out<=159;
				end
				if(in == 3) begin
					state<=5288;
					out<=160;
				end
				if(in == 4) begin
					state<=1399;
					out<=161;
				end
			end
			6074: begin
				if(in == 0) begin
					state<=7221;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=3332;
					out<=164;
				end
				if(in == 3) begin
					state<=5289;
					out<=165;
				end
				if(in == 4) begin
					state<=1400;
					out<=166;
				end
			end
			6075: begin
				if(in == 0) begin
					state<=7212;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=3323;
					out<=169;
				end
				if(in == 3) begin
					state<=5280;
					out<=170;
				end
				if(in == 4) begin
					state<=1391;
					out<=171;
				end
			end
			6076: begin
				if(in == 0) begin
					state<=6087;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=2198;
					out<=174;
				end
				if(in == 3) begin
					state<=4098;
					out<=175;
				end
				if(in == 4) begin
					state<=200;
					out<=176;
				end
			end
			6077: begin
				if(in == 0) begin
					state<=6088;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=2199;
					out<=179;
				end
				if(in == 3) begin
					state<=4099;
					out<=180;
				end
				if(in == 4) begin
					state<=201;
					out<=181;
				end
			end
			6078: begin
				if(in == 0) begin
					state<=6089;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=2200;
					out<=184;
				end
				if(in == 3) begin
					state<=4100;
					out<=185;
				end
				if(in == 4) begin
					state<=202;
					out<=186;
				end
			end
			6079: begin
				if(in == 0) begin
					state<=6090;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=2201;
					out<=189;
				end
				if(in == 3) begin
					state<=4101;
					out<=190;
				end
				if(in == 4) begin
					state<=203;
					out<=191;
				end
			end
			6080: begin
				if(in == 0) begin
					state<=6091;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=2202;
					out<=194;
				end
				if(in == 3) begin
					state<=4102;
					out<=195;
				end
				if(in == 4) begin
					state<=204;
					out<=196;
				end
			end
			6081: begin
				if(in == 0) begin
					state<=6092;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=2203;
					out<=199;
				end
				if(in == 3) begin
					state<=4103;
					out<=200;
				end
				if(in == 4) begin
					state<=205;
					out<=201;
				end
			end
			6082: begin
				if(in == 0) begin
					state<=6093;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=2204;
					out<=204;
				end
				if(in == 3) begin
					state<=4104;
					out<=205;
				end
				if(in == 4) begin
					state<=206;
					out<=206;
				end
			end
			6083: begin
				if(in == 0) begin
					state<=6094;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=2205;
					out<=209;
				end
				if(in == 3) begin
					state<=4105;
					out<=210;
				end
				if(in == 4) begin
					state<=207;
					out<=211;
				end
			end
			6084: begin
				if(in == 0) begin
					state<=6085;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=2196;
					out<=214;
				end
				if(in == 3) begin
					state<=4096;
					out<=215;
				end
				if(in == 4) begin
					state<=198;
					out<=216;
				end
			end
			6085: begin
				if(in == 0) begin
					state<=6096;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=2207;
					out<=219;
				end
				if(in == 3) begin
					state<=4107;
					out<=220;
				end
				if(in == 4) begin
					state<=209;
					out<=221;
				end
			end
			6086: begin
				if(in == 0) begin
					state<=6097;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=2208;
					out<=224;
				end
				if(in == 3) begin
					state<=4108;
					out<=225;
				end
				if(in == 4) begin
					state<=210;
					out<=226;
				end
			end
			6087: begin
				if(in == 0) begin
					state<=6098;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=2209;
					out<=229;
				end
				if(in == 3) begin
					state<=4109;
					out<=230;
				end
				if(in == 4) begin
					state<=211;
					out<=231;
				end
			end
			6088: begin
				if(in == 0) begin
					state<=6099;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=2210;
					out<=234;
				end
				if(in == 3) begin
					state<=4110;
					out<=235;
				end
				if(in == 4) begin
					state<=212;
					out<=236;
				end
			end
			6089: begin
				if(in == 0) begin
					state<=6100;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=2211;
					out<=239;
				end
				if(in == 3) begin
					state<=4111;
					out<=240;
				end
				if(in == 4) begin
					state<=213;
					out<=241;
				end
			end
			6090: begin
				if(in == 0) begin
					state<=6101;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=2212;
					out<=244;
				end
				if(in == 3) begin
					state<=4112;
					out<=245;
				end
				if(in == 4) begin
					state<=214;
					out<=246;
				end
			end
			6091: begin
				if(in == 0) begin
					state<=6102;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=2213;
					out<=249;
				end
				if(in == 3) begin
					state<=4113;
					out<=250;
				end
				if(in == 4) begin
					state<=215;
					out<=251;
				end
			end
			6092: begin
				if(in == 0) begin
					state<=6103;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=2214;
					out<=254;
				end
				if(in == 3) begin
					state<=4114;
					out<=255;
				end
				if(in == 4) begin
					state<=216;
					out<=0;
				end
			end
			6093: begin
				if(in == 0) begin
					state<=6104;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=2215;
					out<=3;
				end
				if(in == 3) begin
					state<=4115;
					out<=4;
				end
				if(in == 4) begin
					state<=217;
					out<=5;
				end
			end
			6094: begin
				if(in == 0) begin
					state<=6095;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=2206;
					out<=8;
				end
				if(in == 3) begin
					state<=4106;
					out<=9;
				end
				if(in == 4) begin
					state<=208;
					out<=10;
				end
			end
			6095: begin
				if(in == 0) begin
					state<=6106;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=2217;
					out<=13;
				end
				if(in == 3) begin
					state<=4117;
					out<=14;
				end
				if(in == 4) begin
					state<=219;
					out<=15;
				end
			end
			6096: begin
				if(in == 0) begin
					state<=6107;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=2218;
					out<=18;
				end
				if(in == 3) begin
					state<=4118;
					out<=19;
				end
				if(in == 4) begin
					state<=220;
					out<=20;
				end
			end
			6097: begin
				if(in == 0) begin
					state<=6108;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=2219;
					out<=23;
				end
				if(in == 3) begin
					state<=4119;
					out<=24;
				end
				if(in == 4) begin
					state<=221;
					out<=25;
				end
			end
			6098: begin
				if(in == 0) begin
					state<=6109;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=2220;
					out<=28;
				end
				if(in == 3) begin
					state<=4120;
					out<=29;
				end
				if(in == 4) begin
					state<=222;
					out<=30;
				end
			end
			6099: begin
				if(in == 0) begin
					state<=6110;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=2221;
					out<=33;
				end
				if(in == 3) begin
					state<=4121;
					out<=34;
				end
				if(in == 4) begin
					state<=223;
					out<=35;
				end
			end
			6100: begin
				if(in == 0) begin
					state<=6111;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=2222;
					out<=38;
				end
				if(in == 3) begin
					state<=4122;
					out<=39;
				end
				if(in == 4) begin
					state<=224;
					out<=40;
				end
			end
			6101: begin
				if(in == 0) begin
					state<=6112;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=2223;
					out<=43;
				end
				if(in == 3) begin
					state<=4123;
					out<=44;
				end
				if(in == 4) begin
					state<=225;
					out<=45;
				end
			end
			6102: begin
				if(in == 0) begin
					state<=6113;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=2224;
					out<=48;
				end
				if(in == 3) begin
					state<=4124;
					out<=49;
				end
				if(in == 4) begin
					state<=226;
					out<=50;
				end
			end
			6103: begin
				if(in == 0) begin
					state<=6114;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=2225;
					out<=53;
				end
				if(in == 3) begin
					state<=4125;
					out<=54;
				end
				if(in == 4) begin
					state<=227;
					out<=55;
				end
			end
			6104: begin
				if(in == 0) begin
					state<=6105;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=2216;
					out<=58;
				end
				if(in == 3) begin
					state<=4116;
					out<=59;
				end
				if(in == 4) begin
					state<=218;
					out<=60;
				end
			end
			6105: begin
				if(in == 0) begin
					state<=6116;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=2227;
					out<=63;
				end
				if(in == 3) begin
					state<=4127;
					out<=64;
				end
				if(in == 4) begin
					state<=229;
					out<=65;
				end
			end
			6106: begin
				if(in == 0) begin
					state<=6117;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=2228;
					out<=68;
				end
				if(in == 3) begin
					state<=4128;
					out<=69;
				end
				if(in == 4) begin
					state<=230;
					out<=70;
				end
			end
			6107: begin
				if(in == 0) begin
					state<=6118;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=2229;
					out<=73;
				end
				if(in == 3) begin
					state<=4129;
					out<=74;
				end
				if(in == 4) begin
					state<=231;
					out<=75;
				end
			end
			6108: begin
				if(in == 0) begin
					state<=6119;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=2230;
					out<=78;
				end
				if(in == 3) begin
					state<=4130;
					out<=79;
				end
				if(in == 4) begin
					state<=232;
					out<=80;
				end
			end
			6109: begin
				if(in == 0) begin
					state<=6120;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=2231;
					out<=83;
				end
				if(in == 3) begin
					state<=4131;
					out<=84;
				end
				if(in == 4) begin
					state<=233;
					out<=85;
				end
			end
			6110: begin
				if(in == 0) begin
					state<=6121;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=2232;
					out<=88;
				end
				if(in == 3) begin
					state<=4132;
					out<=89;
				end
				if(in == 4) begin
					state<=234;
					out<=90;
				end
			end
			6111: begin
				if(in == 0) begin
					state<=6122;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=2233;
					out<=93;
				end
				if(in == 3) begin
					state<=4133;
					out<=94;
				end
				if(in == 4) begin
					state<=235;
					out<=95;
				end
			end
			6112: begin
				if(in == 0) begin
					state<=6123;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=2234;
					out<=98;
				end
				if(in == 3) begin
					state<=4134;
					out<=99;
				end
				if(in == 4) begin
					state<=236;
					out<=100;
				end
			end
			6113: begin
				if(in == 0) begin
					state<=6124;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=2235;
					out<=103;
				end
				if(in == 3) begin
					state<=4135;
					out<=104;
				end
				if(in == 4) begin
					state<=237;
					out<=105;
				end
			end
			6114: begin
				if(in == 0) begin
					state<=6115;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=2226;
					out<=108;
				end
				if(in == 3) begin
					state<=4126;
					out<=109;
				end
				if(in == 4) begin
					state<=228;
					out<=110;
				end
			end
			6115: begin
				if(in == 0) begin
					state<=6126;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=2237;
					out<=113;
				end
				if(in == 3) begin
					state<=4137;
					out<=114;
				end
				if(in == 4) begin
					state<=239;
					out<=115;
				end
			end
			6116: begin
				if(in == 0) begin
					state<=6127;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=2238;
					out<=118;
				end
				if(in == 3) begin
					state<=4138;
					out<=119;
				end
				if(in == 4) begin
					state<=240;
					out<=120;
				end
			end
			6117: begin
				if(in == 0) begin
					state<=6128;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=2239;
					out<=123;
				end
				if(in == 3) begin
					state<=4139;
					out<=124;
				end
				if(in == 4) begin
					state<=241;
					out<=125;
				end
			end
			6118: begin
				if(in == 0) begin
					state<=6129;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=2240;
					out<=128;
				end
				if(in == 3) begin
					state<=4140;
					out<=129;
				end
				if(in == 4) begin
					state<=242;
					out<=130;
				end
			end
			6119: begin
				if(in == 0) begin
					state<=6130;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=2241;
					out<=133;
				end
				if(in == 3) begin
					state<=4141;
					out<=134;
				end
				if(in == 4) begin
					state<=243;
					out<=135;
				end
			end
			6120: begin
				if(in == 0) begin
					state<=6131;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=2242;
					out<=138;
				end
				if(in == 3) begin
					state<=4142;
					out<=139;
				end
				if(in == 4) begin
					state<=244;
					out<=140;
				end
			end
			6121: begin
				if(in == 0) begin
					state<=6132;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=2243;
					out<=143;
				end
				if(in == 3) begin
					state<=4143;
					out<=144;
				end
				if(in == 4) begin
					state<=245;
					out<=145;
				end
			end
			6122: begin
				if(in == 0) begin
					state<=6133;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=2244;
					out<=148;
				end
				if(in == 3) begin
					state<=4144;
					out<=149;
				end
				if(in == 4) begin
					state<=246;
					out<=150;
				end
			end
			6123: begin
				if(in == 0) begin
					state<=6134;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=2245;
					out<=153;
				end
				if(in == 3) begin
					state<=4145;
					out<=154;
				end
				if(in == 4) begin
					state<=247;
					out<=155;
				end
			end
			6124: begin
				if(in == 0) begin
					state<=6125;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=2236;
					out<=158;
				end
				if(in == 3) begin
					state<=4136;
					out<=159;
				end
				if(in == 4) begin
					state<=238;
					out<=160;
				end
			end
			6125: begin
				if(in == 0) begin
					state<=6136;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=2247;
					out<=163;
				end
				if(in == 3) begin
					state<=4147;
					out<=164;
				end
				if(in == 4) begin
					state<=249;
					out<=165;
				end
			end
			6126: begin
				if(in == 0) begin
					state<=6137;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=2248;
					out<=168;
				end
				if(in == 3) begin
					state<=4148;
					out<=169;
				end
				if(in == 4) begin
					state<=250;
					out<=170;
				end
			end
			6127: begin
				if(in == 0) begin
					state<=6138;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=2249;
					out<=173;
				end
				if(in == 3) begin
					state<=4149;
					out<=174;
				end
				if(in == 4) begin
					state<=251;
					out<=175;
				end
			end
			6128: begin
				if(in == 0) begin
					state<=6139;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=2250;
					out<=178;
				end
				if(in == 3) begin
					state<=4150;
					out<=179;
				end
				if(in == 4) begin
					state<=252;
					out<=180;
				end
			end
			6129: begin
				if(in == 0) begin
					state<=6140;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=2251;
					out<=183;
				end
				if(in == 3) begin
					state<=4151;
					out<=184;
				end
				if(in == 4) begin
					state<=253;
					out<=185;
				end
			end
			6130: begin
				if(in == 0) begin
					state<=6141;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=2252;
					out<=188;
				end
				if(in == 3) begin
					state<=4152;
					out<=189;
				end
				if(in == 4) begin
					state<=254;
					out<=190;
				end
			end
			6131: begin
				if(in == 0) begin
					state<=6142;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=2253;
					out<=193;
				end
				if(in == 3) begin
					state<=4153;
					out<=194;
				end
				if(in == 4) begin
					state<=255;
					out<=195;
				end
			end
			6132: begin
				if(in == 0) begin
					state<=6143;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=2254;
					out<=198;
				end
				if(in == 3) begin
					state<=4154;
					out<=199;
				end
				if(in == 4) begin
					state<=256;
					out<=200;
				end
			end
			6133: begin
				if(in == 0) begin
					state<=6144;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=2255;
					out<=203;
				end
				if(in == 3) begin
					state<=4155;
					out<=204;
				end
				if(in == 4) begin
					state<=257;
					out<=205;
				end
			end
			6134: begin
				if(in == 0) begin
					state<=6135;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=2246;
					out<=208;
				end
				if(in == 3) begin
					state<=4146;
					out<=209;
				end
				if(in == 4) begin
					state<=248;
					out<=210;
				end
			end
			6135: begin
				if(in == 0) begin
					state<=7244;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=3355;
					out<=213;
				end
				if(in == 3) begin
					state<=5312;
					out<=214;
				end
				if(in == 4) begin
					state<=1423;
					out<=215;
				end
			end
			6136: begin
				if(in == 0) begin
					state<=7245;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=3356;
					out<=218;
				end
				if(in == 3) begin
					state<=5313;
					out<=219;
				end
				if(in == 4) begin
					state<=1424;
					out<=220;
				end
			end
			6137: begin
				if(in == 0) begin
					state<=7246;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=3357;
					out<=223;
				end
				if(in == 3) begin
					state<=5314;
					out<=224;
				end
				if(in == 4) begin
					state<=1425;
					out<=225;
				end
			end
			6138: begin
				if(in == 0) begin
					state<=7247;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=3358;
					out<=228;
				end
				if(in == 3) begin
					state<=5315;
					out<=229;
				end
				if(in == 4) begin
					state<=1426;
					out<=230;
				end
			end
			6139: begin
				if(in == 0) begin
					state<=7248;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=3359;
					out<=233;
				end
				if(in == 3) begin
					state<=5316;
					out<=234;
				end
				if(in == 4) begin
					state<=1427;
					out<=235;
				end
			end
			6140: begin
				if(in == 0) begin
					state<=7249;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=3360;
					out<=238;
				end
				if(in == 3) begin
					state<=5317;
					out<=239;
				end
				if(in == 4) begin
					state<=1428;
					out<=240;
				end
			end
			6141: begin
				if(in == 0) begin
					state<=7250;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=3361;
					out<=243;
				end
				if(in == 3) begin
					state<=5318;
					out<=244;
				end
				if(in == 4) begin
					state<=1429;
					out<=245;
				end
			end
			6142: begin
				if(in == 0) begin
					state<=7251;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=3362;
					out<=248;
				end
				if(in == 3) begin
					state<=5319;
					out<=249;
				end
				if(in == 4) begin
					state<=1430;
					out<=250;
				end
			end
			6143: begin
				if(in == 0) begin
					state<=7252;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=3363;
					out<=253;
				end
				if(in == 3) begin
					state<=5320;
					out<=254;
				end
				if(in == 4) begin
					state<=1431;
					out<=255;
				end
			end
			6144: begin
				if(in == 0) begin
					state<=7243;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=3354;
					out<=2;
				end
				if(in == 3) begin
					state<=5311;
					out<=3;
				end
				if(in == 4) begin
					state<=1422;
					out<=4;
				end
			end
			6145: begin
				if(in == 0) begin
					state<=6156;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=2267;
					out<=7;
				end
				if(in == 3) begin
					state<=4167;
					out<=8;
				end
				if(in == 4) begin
					state<=269;
					out<=9;
				end
			end
			6146: begin
				if(in == 0) begin
					state<=6157;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=2268;
					out<=12;
				end
				if(in == 3) begin
					state<=4168;
					out<=13;
				end
				if(in == 4) begin
					state<=270;
					out<=14;
				end
			end
			6147: begin
				if(in == 0) begin
					state<=6158;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=2269;
					out<=17;
				end
				if(in == 3) begin
					state<=4169;
					out<=18;
				end
				if(in == 4) begin
					state<=271;
					out<=19;
				end
			end
			6148: begin
				if(in == 0) begin
					state<=6159;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=2270;
					out<=22;
				end
				if(in == 3) begin
					state<=4170;
					out<=23;
				end
				if(in == 4) begin
					state<=272;
					out<=24;
				end
			end
			6149: begin
				if(in == 0) begin
					state<=6160;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=2271;
					out<=27;
				end
				if(in == 3) begin
					state<=4171;
					out<=28;
				end
				if(in == 4) begin
					state<=273;
					out<=29;
				end
			end
			6150: begin
				if(in == 0) begin
					state<=6161;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=2272;
					out<=32;
				end
				if(in == 3) begin
					state<=4172;
					out<=33;
				end
				if(in == 4) begin
					state<=274;
					out<=34;
				end
			end
			6151: begin
				if(in == 0) begin
					state<=6162;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=2273;
					out<=37;
				end
				if(in == 3) begin
					state<=4173;
					out<=38;
				end
				if(in == 4) begin
					state<=275;
					out<=39;
				end
			end
			6152: begin
				if(in == 0) begin
					state<=6163;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=2274;
					out<=42;
				end
				if(in == 3) begin
					state<=4174;
					out<=43;
				end
				if(in == 4) begin
					state<=276;
					out<=44;
				end
			end
			6153: begin
				if(in == 0) begin
					state<=6154;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=2265;
					out<=47;
				end
				if(in == 3) begin
					state<=4165;
					out<=48;
				end
				if(in == 4) begin
					state<=267;
					out<=49;
				end
			end
			6154: begin
				if(in == 0) begin
					state<=6165;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=2276;
					out<=52;
				end
				if(in == 3) begin
					state<=4176;
					out<=53;
				end
				if(in == 4) begin
					state<=278;
					out<=54;
				end
			end
			6155: begin
				if(in == 0) begin
					state<=6166;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=2277;
					out<=57;
				end
				if(in == 3) begin
					state<=4177;
					out<=58;
				end
				if(in == 4) begin
					state<=279;
					out<=59;
				end
			end
			6156: begin
				if(in == 0) begin
					state<=6167;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=2278;
					out<=62;
				end
				if(in == 3) begin
					state<=4178;
					out<=63;
				end
				if(in == 4) begin
					state<=280;
					out<=64;
				end
			end
			6157: begin
				if(in == 0) begin
					state<=6168;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=2279;
					out<=67;
				end
				if(in == 3) begin
					state<=4179;
					out<=68;
				end
				if(in == 4) begin
					state<=281;
					out<=69;
				end
			end
			6158: begin
				if(in == 0) begin
					state<=6169;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=2280;
					out<=72;
				end
				if(in == 3) begin
					state<=4180;
					out<=73;
				end
				if(in == 4) begin
					state<=282;
					out<=74;
				end
			end
			6159: begin
				if(in == 0) begin
					state<=6170;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=2281;
					out<=77;
				end
				if(in == 3) begin
					state<=4181;
					out<=78;
				end
				if(in == 4) begin
					state<=283;
					out<=79;
				end
			end
			6160: begin
				if(in == 0) begin
					state<=6171;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=2282;
					out<=82;
				end
				if(in == 3) begin
					state<=4182;
					out<=83;
				end
				if(in == 4) begin
					state<=284;
					out<=84;
				end
			end
			6161: begin
				if(in == 0) begin
					state<=6172;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=2283;
					out<=87;
				end
				if(in == 3) begin
					state<=4183;
					out<=88;
				end
				if(in == 4) begin
					state<=285;
					out<=89;
				end
			end
			6162: begin
				if(in == 0) begin
					state<=6173;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=2284;
					out<=92;
				end
				if(in == 3) begin
					state<=4184;
					out<=93;
				end
				if(in == 4) begin
					state<=286;
					out<=94;
				end
			end
			6163: begin
				if(in == 0) begin
					state<=6164;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=2275;
					out<=97;
				end
				if(in == 3) begin
					state<=4175;
					out<=98;
				end
				if(in == 4) begin
					state<=277;
					out<=99;
				end
			end
			6164: begin
				if(in == 0) begin
					state<=6175;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=2286;
					out<=102;
				end
				if(in == 3) begin
					state<=4186;
					out<=103;
				end
				if(in == 4) begin
					state<=288;
					out<=104;
				end
			end
			6165: begin
				if(in == 0) begin
					state<=6176;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=2287;
					out<=107;
				end
				if(in == 3) begin
					state<=4187;
					out<=108;
				end
				if(in == 4) begin
					state<=289;
					out<=109;
				end
			end
			6166: begin
				if(in == 0) begin
					state<=6177;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=2288;
					out<=112;
				end
				if(in == 3) begin
					state<=4188;
					out<=113;
				end
				if(in == 4) begin
					state<=290;
					out<=114;
				end
			end
			6167: begin
				if(in == 0) begin
					state<=6178;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=2289;
					out<=117;
				end
				if(in == 3) begin
					state<=4189;
					out<=118;
				end
				if(in == 4) begin
					state<=291;
					out<=119;
				end
			end
			6168: begin
				if(in == 0) begin
					state<=6179;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=2290;
					out<=122;
				end
				if(in == 3) begin
					state<=4190;
					out<=123;
				end
				if(in == 4) begin
					state<=292;
					out<=124;
				end
			end
			6169: begin
				if(in == 0) begin
					state<=6180;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=2291;
					out<=127;
				end
				if(in == 3) begin
					state<=4191;
					out<=128;
				end
				if(in == 4) begin
					state<=293;
					out<=129;
				end
			end
			6170: begin
				if(in == 0) begin
					state<=6181;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=2292;
					out<=132;
				end
				if(in == 3) begin
					state<=4192;
					out<=133;
				end
				if(in == 4) begin
					state<=294;
					out<=134;
				end
			end
			6171: begin
				if(in == 0) begin
					state<=6182;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=2293;
					out<=137;
				end
				if(in == 3) begin
					state<=4193;
					out<=138;
				end
				if(in == 4) begin
					state<=295;
					out<=139;
				end
			end
			6172: begin
				if(in == 0) begin
					state<=6183;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=2294;
					out<=142;
				end
				if(in == 3) begin
					state<=4194;
					out<=143;
				end
				if(in == 4) begin
					state<=296;
					out<=144;
				end
			end
			6173: begin
				if(in == 0) begin
					state<=6174;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=2285;
					out<=147;
				end
				if(in == 3) begin
					state<=4185;
					out<=148;
				end
				if(in == 4) begin
					state<=287;
					out<=149;
				end
			end
			6174: begin
				if(in == 0) begin
					state<=6185;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=2296;
					out<=152;
				end
				if(in == 3) begin
					state<=4196;
					out<=153;
				end
				if(in == 4) begin
					state<=298;
					out<=154;
				end
			end
			6175: begin
				if(in == 0) begin
					state<=6186;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=2297;
					out<=157;
				end
				if(in == 3) begin
					state<=4197;
					out<=158;
				end
				if(in == 4) begin
					state<=299;
					out<=159;
				end
			end
			6176: begin
				if(in == 0) begin
					state<=6187;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=2298;
					out<=162;
				end
				if(in == 3) begin
					state<=4198;
					out<=163;
				end
				if(in == 4) begin
					state<=300;
					out<=164;
				end
			end
			6177: begin
				if(in == 0) begin
					state<=6188;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=2299;
					out<=167;
				end
				if(in == 3) begin
					state<=4199;
					out<=168;
				end
				if(in == 4) begin
					state<=301;
					out<=169;
				end
			end
			6178: begin
				if(in == 0) begin
					state<=6189;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=2300;
					out<=172;
				end
				if(in == 3) begin
					state<=4200;
					out<=173;
				end
				if(in == 4) begin
					state<=302;
					out<=174;
				end
			end
			6179: begin
				if(in == 0) begin
					state<=6190;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=2301;
					out<=177;
				end
				if(in == 3) begin
					state<=4201;
					out<=178;
				end
				if(in == 4) begin
					state<=303;
					out<=179;
				end
			end
			6180: begin
				if(in == 0) begin
					state<=6191;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=2302;
					out<=182;
				end
				if(in == 3) begin
					state<=4202;
					out<=183;
				end
				if(in == 4) begin
					state<=304;
					out<=184;
				end
			end
			6181: begin
				if(in == 0) begin
					state<=6192;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=2303;
					out<=187;
				end
				if(in == 3) begin
					state<=4203;
					out<=188;
				end
				if(in == 4) begin
					state<=305;
					out<=189;
				end
			end
			6182: begin
				if(in == 0) begin
					state<=6193;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=2304;
					out<=192;
				end
				if(in == 3) begin
					state<=4204;
					out<=193;
				end
				if(in == 4) begin
					state<=306;
					out<=194;
				end
			end
			6183: begin
				if(in == 0) begin
					state<=6184;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=2295;
					out<=197;
				end
				if(in == 3) begin
					state<=4195;
					out<=198;
				end
				if(in == 4) begin
					state<=297;
					out<=199;
				end
			end
			6184: begin
				if(in == 0) begin
					state<=6195;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=2306;
					out<=202;
				end
				if(in == 3) begin
					state<=4206;
					out<=203;
				end
				if(in == 4) begin
					state<=308;
					out<=204;
				end
			end
			6185: begin
				if(in == 0) begin
					state<=6196;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=2307;
					out<=207;
				end
				if(in == 3) begin
					state<=4207;
					out<=208;
				end
				if(in == 4) begin
					state<=309;
					out<=209;
				end
			end
			6186: begin
				if(in == 0) begin
					state<=6197;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=2308;
					out<=212;
				end
				if(in == 3) begin
					state<=4208;
					out<=213;
				end
				if(in == 4) begin
					state<=310;
					out<=214;
				end
			end
			6187: begin
				if(in == 0) begin
					state<=6198;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=2309;
					out<=217;
				end
				if(in == 3) begin
					state<=4209;
					out<=218;
				end
				if(in == 4) begin
					state<=311;
					out<=219;
				end
			end
			6188: begin
				if(in == 0) begin
					state<=6199;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=2310;
					out<=222;
				end
				if(in == 3) begin
					state<=4210;
					out<=223;
				end
				if(in == 4) begin
					state<=312;
					out<=224;
				end
			end
			6189: begin
				if(in == 0) begin
					state<=6200;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=2311;
					out<=227;
				end
				if(in == 3) begin
					state<=4211;
					out<=228;
				end
				if(in == 4) begin
					state<=313;
					out<=229;
				end
			end
			6190: begin
				if(in == 0) begin
					state<=6201;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=2312;
					out<=232;
				end
				if(in == 3) begin
					state<=4212;
					out<=233;
				end
				if(in == 4) begin
					state<=314;
					out<=234;
				end
			end
			6191: begin
				if(in == 0) begin
					state<=6202;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=2313;
					out<=237;
				end
				if(in == 3) begin
					state<=4213;
					out<=238;
				end
				if(in == 4) begin
					state<=315;
					out<=239;
				end
			end
			6192: begin
				if(in == 0) begin
					state<=6203;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=2314;
					out<=242;
				end
				if(in == 3) begin
					state<=4214;
					out<=243;
				end
				if(in == 4) begin
					state<=316;
					out<=244;
				end
			end
			6193: begin
				if(in == 0) begin
					state<=6194;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=2305;
					out<=247;
				end
				if(in == 3) begin
					state<=4205;
					out<=248;
				end
				if(in == 4) begin
					state<=307;
					out<=249;
				end
			end
			6194: begin
				if(in == 0) begin
					state<=6205;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=2316;
					out<=252;
				end
				if(in == 3) begin
					state<=4216;
					out<=253;
				end
				if(in == 4) begin
					state<=318;
					out<=254;
				end
			end
			6195: begin
				if(in == 0) begin
					state<=6206;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=2317;
					out<=1;
				end
				if(in == 3) begin
					state<=4217;
					out<=2;
				end
				if(in == 4) begin
					state<=319;
					out<=3;
				end
			end
			6196: begin
				if(in == 0) begin
					state<=6207;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=2318;
					out<=6;
				end
				if(in == 3) begin
					state<=4218;
					out<=7;
				end
				if(in == 4) begin
					state<=320;
					out<=8;
				end
			end
			6197: begin
				if(in == 0) begin
					state<=6208;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=2319;
					out<=11;
				end
				if(in == 3) begin
					state<=4219;
					out<=12;
				end
				if(in == 4) begin
					state<=321;
					out<=13;
				end
			end
			6198: begin
				if(in == 0) begin
					state<=6209;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=2320;
					out<=16;
				end
				if(in == 3) begin
					state<=4220;
					out<=17;
				end
				if(in == 4) begin
					state<=322;
					out<=18;
				end
			end
			6199: begin
				if(in == 0) begin
					state<=6210;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=2321;
					out<=21;
				end
				if(in == 3) begin
					state<=4221;
					out<=22;
				end
				if(in == 4) begin
					state<=323;
					out<=23;
				end
			end
			6200: begin
				if(in == 0) begin
					state<=6211;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=2322;
					out<=26;
				end
				if(in == 3) begin
					state<=4222;
					out<=27;
				end
				if(in == 4) begin
					state<=324;
					out<=28;
				end
			end
			6201: begin
				if(in == 0) begin
					state<=6212;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=2323;
					out<=31;
				end
				if(in == 3) begin
					state<=4223;
					out<=32;
				end
				if(in == 4) begin
					state<=325;
					out<=33;
				end
			end
			6202: begin
				if(in == 0) begin
					state<=6213;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=2324;
					out<=36;
				end
				if(in == 3) begin
					state<=4224;
					out<=37;
				end
				if(in == 4) begin
					state<=326;
					out<=38;
				end
			end
			6203: begin
				if(in == 0) begin
					state<=6204;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=2315;
					out<=41;
				end
				if(in == 3) begin
					state<=4215;
					out<=42;
				end
				if(in == 4) begin
					state<=317;
					out<=43;
				end
			end
			6204: begin
				if(in == 0) begin
					state<=6788;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=2899;
					out<=46;
				end
				if(in == 3) begin
					state<=5343;
					out<=47;
				end
				if(in == 4) begin
					state<=1454;
					out<=48;
				end
			end
			6205: begin
				if(in == 0) begin
					state<=6789;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=2900;
					out<=51;
				end
				if(in == 3) begin
					state<=5344;
					out<=52;
				end
				if(in == 4) begin
					state<=1455;
					out<=53;
				end
			end
			6206: begin
				if(in == 0) begin
					state<=6790;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=2901;
					out<=56;
				end
				if(in == 3) begin
					state<=5345;
					out<=57;
				end
				if(in == 4) begin
					state<=1456;
					out<=58;
				end
			end
			6207: begin
				if(in == 0) begin
					state<=6791;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=2902;
					out<=61;
				end
				if(in == 3) begin
					state<=5346;
					out<=62;
				end
				if(in == 4) begin
					state<=1457;
					out<=63;
				end
			end
			6208: begin
				if(in == 0) begin
					state<=6792;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=2903;
					out<=66;
				end
				if(in == 3) begin
					state<=5347;
					out<=67;
				end
				if(in == 4) begin
					state<=1458;
					out<=68;
				end
			end
			6209: begin
				if(in == 0) begin
					state<=6793;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=2904;
					out<=71;
				end
				if(in == 3) begin
					state<=5348;
					out<=72;
				end
				if(in == 4) begin
					state<=1459;
					out<=73;
				end
			end
			6210: begin
				if(in == 0) begin
					state<=6794;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=2905;
					out<=76;
				end
				if(in == 3) begin
					state<=5349;
					out<=77;
				end
				if(in == 4) begin
					state<=1460;
					out<=78;
				end
			end
			6211: begin
				if(in == 0) begin
					state<=6795;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=2906;
					out<=81;
				end
				if(in == 3) begin
					state<=5350;
					out<=82;
				end
				if(in == 4) begin
					state<=1461;
					out<=83;
				end
			end
			6212: begin
				if(in == 0) begin
					state<=6796;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=2907;
					out<=86;
				end
				if(in == 3) begin
					state<=5351;
					out<=87;
				end
				if(in == 4) begin
					state<=1462;
					out<=88;
				end
			end
			6213: begin
				if(in == 0) begin
					state<=6787;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=2898;
					out<=91;
				end
				if(in == 3) begin
					state<=5342;
					out<=92;
				end
				if(in == 4) begin
					state<=1453;
					out<=93;
				end
			end
			6214: begin
				if(in == 0) begin
					state<=6225;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=2336;
					out<=96;
				end
				if(in == 3) begin
					state<=4236;
					out<=97;
				end
				if(in == 4) begin
					state<=338;
					out<=98;
				end
			end
			6215: begin
				if(in == 0) begin
					state<=6226;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=2337;
					out<=101;
				end
				if(in == 3) begin
					state<=4237;
					out<=102;
				end
				if(in == 4) begin
					state<=339;
					out<=103;
				end
			end
			6216: begin
				if(in == 0) begin
					state<=6227;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=2338;
					out<=106;
				end
				if(in == 3) begin
					state<=4238;
					out<=107;
				end
				if(in == 4) begin
					state<=340;
					out<=108;
				end
			end
			6217: begin
				if(in == 0) begin
					state<=6228;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=2339;
					out<=111;
				end
				if(in == 3) begin
					state<=4239;
					out<=112;
				end
				if(in == 4) begin
					state<=341;
					out<=113;
				end
			end
			6218: begin
				if(in == 0) begin
					state<=6229;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=2340;
					out<=116;
				end
				if(in == 3) begin
					state<=4240;
					out<=117;
				end
				if(in == 4) begin
					state<=342;
					out<=118;
				end
			end
			6219: begin
				if(in == 0) begin
					state<=6230;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=2341;
					out<=121;
				end
				if(in == 3) begin
					state<=4241;
					out<=122;
				end
				if(in == 4) begin
					state<=343;
					out<=123;
				end
			end
			6220: begin
				if(in == 0) begin
					state<=6231;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=2342;
					out<=126;
				end
				if(in == 3) begin
					state<=4242;
					out<=127;
				end
				if(in == 4) begin
					state<=344;
					out<=128;
				end
			end
			6221: begin
				if(in == 0) begin
					state<=6232;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=2343;
					out<=131;
				end
				if(in == 3) begin
					state<=4243;
					out<=132;
				end
				if(in == 4) begin
					state<=345;
					out<=133;
				end
			end
			6222: begin
				if(in == 0) begin
					state<=6223;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=2334;
					out<=136;
				end
				if(in == 3) begin
					state<=4234;
					out<=137;
				end
				if(in == 4) begin
					state<=336;
					out<=138;
				end
			end
			6223: begin
				if(in == 0) begin
					state<=6234;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=2345;
					out<=141;
				end
				if(in == 3) begin
					state<=4245;
					out<=142;
				end
				if(in == 4) begin
					state<=347;
					out<=143;
				end
			end
			6224: begin
				if(in == 0) begin
					state<=6235;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=2346;
					out<=146;
				end
				if(in == 3) begin
					state<=4246;
					out<=147;
				end
				if(in == 4) begin
					state<=348;
					out<=148;
				end
			end
			6225: begin
				if(in == 0) begin
					state<=6236;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=2347;
					out<=151;
				end
				if(in == 3) begin
					state<=4247;
					out<=152;
				end
				if(in == 4) begin
					state<=349;
					out<=153;
				end
			end
			6226: begin
				if(in == 0) begin
					state<=6237;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=2348;
					out<=156;
				end
				if(in == 3) begin
					state<=4248;
					out<=157;
				end
				if(in == 4) begin
					state<=350;
					out<=158;
				end
			end
			6227: begin
				if(in == 0) begin
					state<=6238;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=2349;
					out<=161;
				end
				if(in == 3) begin
					state<=4249;
					out<=162;
				end
				if(in == 4) begin
					state<=351;
					out<=163;
				end
			end
			6228: begin
				if(in == 0) begin
					state<=6239;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=2350;
					out<=166;
				end
				if(in == 3) begin
					state<=4250;
					out<=167;
				end
				if(in == 4) begin
					state<=352;
					out<=168;
				end
			end
			6229: begin
				if(in == 0) begin
					state<=6240;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=2351;
					out<=171;
				end
				if(in == 3) begin
					state<=4251;
					out<=172;
				end
				if(in == 4) begin
					state<=353;
					out<=173;
				end
			end
			6230: begin
				if(in == 0) begin
					state<=6241;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=2352;
					out<=176;
				end
				if(in == 3) begin
					state<=4252;
					out<=177;
				end
				if(in == 4) begin
					state<=354;
					out<=178;
				end
			end
			6231: begin
				if(in == 0) begin
					state<=6242;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=2353;
					out<=181;
				end
				if(in == 3) begin
					state<=4253;
					out<=182;
				end
				if(in == 4) begin
					state<=355;
					out<=183;
				end
			end
			6232: begin
				if(in == 0) begin
					state<=6233;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=2344;
					out<=186;
				end
				if(in == 3) begin
					state<=4244;
					out<=187;
				end
				if(in == 4) begin
					state<=346;
					out<=188;
				end
			end
			6233: begin
				if(in == 0) begin
					state<=6244;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=2355;
					out<=191;
				end
				if(in == 3) begin
					state<=4255;
					out<=192;
				end
				if(in == 4) begin
					state<=357;
					out<=193;
				end
			end
			6234: begin
				if(in == 0) begin
					state<=6245;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=2356;
					out<=196;
				end
				if(in == 3) begin
					state<=4256;
					out<=197;
				end
				if(in == 4) begin
					state<=358;
					out<=198;
				end
			end
			6235: begin
				if(in == 0) begin
					state<=6246;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=2357;
					out<=201;
				end
				if(in == 3) begin
					state<=4257;
					out<=202;
				end
				if(in == 4) begin
					state<=359;
					out<=203;
				end
			end
			6236: begin
				if(in == 0) begin
					state<=6247;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=2358;
					out<=206;
				end
				if(in == 3) begin
					state<=4258;
					out<=207;
				end
				if(in == 4) begin
					state<=360;
					out<=208;
				end
			end
			6237: begin
				if(in == 0) begin
					state<=6248;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=2359;
					out<=211;
				end
				if(in == 3) begin
					state<=4259;
					out<=212;
				end
				if(in == 4) begin
					state<=361;
					out<=213;
				end
			end
			6238: begin
				if(in == 0) begin
					state<=6249;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=2360;
					out<=216;
				end
				if(in == 3) begin
					state<=4260;
					out<=217;
				end
				if(in == 4) begin
					state<=362;
					out<=218;
				end
			end
			6239: begin
				if(in == 0) begin
					state<=6250;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=2361;
					out<=221;
				end
				if(in == 3) begin
					state<=4261;
					out<=222;
				end
				if(in == 4) begin
					state<=363;
					out<=223;
				end
			end
			6240: begin
				if(in == 0) begin
					state<=6251;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=2362;
					out<=226;
				end
				if(in == 3) begin
					state<=4262;
					out<=227;
				end
				if(in == 4) begin
					state<=364;
					out<=228;
				end
			end
			6241: begin
				if(in == 0) begin
					state<=6252;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=2363;
					out<=231;
				end
				if(in == 3) begin
					state<=4263;
					out<=232;
				end
				if(in == 4) begin
					state<=365;
					out<=233;
				end
			end
			6242: begin
				if(in == 0) begin
					state<=6243;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=2354;
					out<=236;
				end
				if(in == 3) begin
					state<=4254;
					out<=237;
				end
				if(in == 4) begin
					state<=356;
					out<=238;
				end
			end
			6243: begin
				if(in == 0) begin
					state<=6254;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=2365;
					out<=241;
				end
				if(in == 3) begin
					state<=4265;
					out<=242;
				end
				if(in == 4) begin
					state<=367;
					out<=243;
				end
			end
			6244: begin
				if(in == 0) begin
					state<=6255;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=2366;
					out<=246;
				end
				if(in == 3) begin
					state<=4266;
					out<=247;
				end
				if(in == 4) begin
					state<=368;
					out<=248;
				end
			end
			6245: begin
				if(in == 0) begin
					state<=6256;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=2367;
					out<=251;
				end
				if(in == 3) begin
					state<=4267;
					out<=252;
				end
				if(in == 4) begin
					state<=369;
					out<=253;
				end
			end
			6246: begin
				if(in == 0) begin
					state<=6257;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=2368;
					out<=0;
				end
				if(in == 3) begin
					state<=4268;
					out<=1;
				end
				if(in == 4) begin
					state<=370;
					out<=2;
				end
			end
			6247: begin
				if(in == 0) begin
					state<=6258;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=2369;
					out<=5;
				end
				if(in == 3) begin
					state<=4269;
					out<=6;
				end
				if(in == 4) begin
					state<=371;
					out<=7;
				end
			end
			6248: begin
				if(in == 0) begin
					state<=6259;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=2370;
					out<=10;
				end
				if(in == 3) begin
					state<=4270;
					out<=11;
				end
				if(in == 4) begin
					state<=372;
					out<=12;
				end
			end
			6249: begin
				if(in == 0) begin
					state<=6260;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=2371;
					out<=15;
				end
				if(in == 3) begin
					state<=4271;
					out<=16;
				end
				if(in == 4) begin
					state<=373;
					out<=17;
				end
			end
			6250: begin
				if(in == 0) begin
					state<=6261;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=2372;
					out<=20;
				end
				if(in == 3) begin
					state<=4272;
					out<=21;
				end
				if(in == 4) begin
					state<=374;
					out<=22;
				end
			end
			6251: begin
				if(in == 0) begin
					state<=6262;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=2373;
					out<=25;
				end
				if(in == 3) begin
					state<=4273;
					out<=26;
				end
				if(in == 4) begin
					state<=375;
					out<=27;
				end
			end
			6252: begin
				if(in == 0) begin
					state<=6253;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=2364;
					out<=30;
				end
				if(in == 3) begin
					state<=4264;
					out<=31;
				end
				if(in == 4) begin
					state<=366;
					out<=32;
				end
			end
			6253: begin
				if(in == 0) begin
					state<=6264;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=2375;
					out<=35;
				end
				if(in == 3) begin
					state<=4275;
					out<=36;
				end
				if(in == 4) begin
					state<=377;
					out<=37;
				end
			end
			6254: begin
				if(in == 0) begin
					state<=6265;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=2376;
					out<=40;
				end
				if(in == 3) begin
					state<=4276;
					out<=41;
				end
				if(in == 4) begin
					state<=378;
					out<=42;
				end
			end
			6255: begin
				if(in == 0) begin
					state<=6266;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=2377;
					out<=45;
				end
				if(in == 3) begin
					state<=4277;
					out<=46;
				end
				if(in == 4) begin
					state<=379;
					out<=47;
				end
			end
			6256: begin
				if(in == 0) begin
					state<=6267;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=2378;
					out<=50;
				end
				if(in == 3) begin
					state<=4278;
					out<=51;
				end
				if(in == 4) begin
					state<=380;
					out<=52;
				end
			end
			6257: begin
				if(in == 0) begin
					state<=6268;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=2379;
					out<=55;
				end
				if(in == 3) begin
					state<=4279;
					out<=56;
				end
				if(in == 4) begin
					state<=381;
					out<=57;
				end
			end
			6258: begin
				if(in == 0) begin
					state<=6269;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=2380;
					out<=60;
				end
				if(in == 3) begin
					state<=4280;
					out<=61;
				end
				if(in == 4) begin
					state<=382;
					out<=62;
				end
			end
			6259: begin
				if(in == 0) begin
					state<=6270;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=2381;
					out<=65;
				end
				if(in == 3) begin
					state<=4281;
					out<=66;
				end
				if(in == 4) begin
					state<=383;
					out<=67;
				end
			end
			6260: begin
				if(in == 0) begin
					state<=6271;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=2382;
					out<=70;
				end
				if(in == 3) begin
					state<=4282;
					out<=71;
				end
				if(in == 4) begin
					state<=384;
					out<=72;
				end
			end
			6261: begin
				if(in == 0) begin
					state<=6272;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=2383;
					out<=75;
				end
				if(in == 3) begin
					state<=4283;
					out<=76;
				end
				if(in == 4) begin
					state<=385;
					out<=77;
				end
			end
			6262: begin
				if(in == 0) begin
					state<=6263;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=2374;
					out<=80;
				end
				if(in == 3) begin
					state<=4274;
					out<=81;
				end
				if(in == 4) begin
					state<=376;
					out<=82;
				end
			end
			6263: begin
				if(in == 0) begin
					state<=6274;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=2385;
					out<=85;
				end
				if(in == 3) begin
					state<=4285;
					out<=86;
				end
				if(in == 4) begin
					state<=387;
					out<=87;
				end
			end
			6264: begin
				if(in == 0) begin
					state<=6275;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=2386;
					out<=90;
				end
				if(in == 3) begin
					state<=4286;
					out<=91;
				end
				if(in == 4) begin
					state<=388;
					out<=92;
				end
			end
			6265: begin
				if(in == 0) begin
					state<=6276;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=2387;
					out<=95;
				end
				if(in == 3) begin
					state<=4287;
					out<=96;
				end
				if(in == 4) begin
					state<=389;
					out<=97;
				end
			end
			6266: begin
				if(in == 0) begin
					state<=6277;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=2388;
					out<=100;
				end
				if(in == 3) begin
					state<=4288;
					out<=101;
				end
				if(in == 4) begin
					state<=390;
					out<=102;
				end
			end
			6267: begin
				if(in == 0) begin
					state<=6278;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=2389;
					out<=105;
				end
				if(in == 3) begin
					state<=4289;
					out<=106;
				end
				if(in == 4) begin
					state<=391;
					out<=107;
				end
			end
			6268: begin
				if(in == 0) begin
					state<=6279;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=2390;
					out<=110;
				end
				if(in == 3) begin
					state<=4290;
					out<=111;
				end
				if(in == 4) begin
					state<=392;
					out<=112;
				end
			end
			6269: begin
				if(in == 0) begin
					state<=6280;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=2391;
					out<=115;
				end
				if(in == 3) begin
					state<=4291;
					out<=116;
				end
				if(in == 4) begin
					state<=393;
					out<=117;
				end
			end
			6270: begin
				if(in == 0) begin
					state<=6281;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=2392;
					out<=120;
				end
				if(in == 3) begin
					state<=4292;
					out<=121;
				end
				if(in == 4) begin
					state<=394;
					out<=122;
				end
			end
			6271: begin
				if(in == 0) begin
					state<=6282;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=2393;
					out<=125;
				end
				if(in == 3) begin
					state<=4293;
					out<=126;
				end
				if(in == 4) begin
					state<=395;
					out<=127;
				end
			end
			6272: begin
				if(in == 0) begin
					state<=6273;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=2384;
					out<=130;
				end
				if(in == 3) begin
					state<=4284;
					out<=131;
				end
				if(in == 4) begin
					state<=386;
					out<=132;
				end
			end
			6273: begin
				if(in == 0) begin
					state<=7275;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=3386;
					out<=135;
				end
				if(in == 3) begin
					state<=4898;
					out<=136;
				end
				if(in == 4) begin
					state<=1000;
					out<=137;
				end
			end
			6274: begin
				if(in == 0) begin
					state<=7276;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=3387;
					out<=140;
				end
				if(in == 3) begin
					state<=4899;
					out<=141;
				end
				if(in == 4) begin
					state<=1001;
					out<=142;
				end
			end
			6275: begin
				if(in == 0) begin
					state<=7277;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=3388;
					out<=145;
				end
				if(in == 3) begin
					state<=4900;
					out<=146;
				end
				if(in == 4) begin
					state<=1002;
					out<=147;
				end
			end
			6276: begin
				if(in == 0) begin
					state<=7278;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=3389;
					out<=150;
				end
				if(in == 3) begin
					state<=4901;
					out<=151;
				end
				if(in == 4) begin
					state<=1003;
					out<=152;
				end
			end
			6277: begin
				if(in == 0) begin
					state<=7279;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=3390;
					out<=155;
				end
				if(in == 3) begin
					state<=4902;
					out<=156;
				end
				if(in == 4) begin
					state<=1004;
					out<=157;
				end
			end
			6278: begin
				if(in == 0) begin
					state<=7280;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=3391;
					out<=160;
				end
				if(in == 3) begin
					state<=4903;
					out<=161;
				end
				if(in == 4) begin
					state<=1005;
					out<=162;
				end
			end
			6279: begin
				if(in == 0) begin
					state<=7281;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=3392;
					out<=165;
				end
				if(in == 3) begin
					state<=4904;
					out<=166;
				end
				if(in == 4) begin
					state<=1006;
					out<=167;
				end
			end
			6280: begin
				if(in == 0) begin
					state<=7282;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=3393;
					out<=170;
				end
				if(in == 3) begin
					state<=4905;
					out<=171;
				end
				if(in == 4) begin
					state<=1007;
					out<=172;
				end
			end
			6281: begin
				if(in == 0) begin
					state<=7283;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=3394;
					out<=175;
				end
				if(in == 3) begin
					state<=4906;
					out<=176;
				end
				if(in == 4) begin
					state<=1008;
					out<=177;
				end
			end
			6282: begin
				if(in == 0) begin
					state<=7274;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=3385;
					out<=180;
				end
				if(in == 3) begin
					state<=4897;
					out<=181;
				end
				if(in == 4) begin
					state<=999;
					out<=182;
				end
			end
			6283: begin
				if(in == 0) begin
					state<=6294;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=2405;
					out<=185;
				end
				if(in == 3) begin
					state<=4305;
					out<=186;
				end
				if(in == 4) begin
					state<=407;
					out<=187;
				end
			end
			6284: begin
				if(in == 0) begin
					state<=6295;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=2406;
					out<=190;
				end
				if(in == 3) begin
					state<=4306;
					out<=191;
				end
				if(in == 4) begin
					state<=408;
					out<=192;
				end
			end
			6285: begin
				if(in == 0) begin
					state<=6296;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=2407;
					out<=195;
				end
				if(in == 3) begin
					state<=4307;
					out<=196;
				end
				if(in == 4) begin
					state<=409;
					out<=197;
				end
			end
			6286: begin
				if(in == 0) begin
					state<=6297;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=2408;
					out<=200;
				end
				if(in == 3) begin
					state<=4308;
					out<=201;
				end
				if(in == 4) begin
					state<=410;
					out<=202;
				end
			end
			6287: begin
				if(in == 0) begin
					state<=6298;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=2409;
					out<=205;
				end
				if(in == 3) begin
					state<=4309;
					out<=206;
				end
				if(in == 4) begin
					state<=411;
					out<=207;
				end
			end
			6288: begin
				if(in == 0) begin
					state<=6299;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=2410;
					out<=210;
				end
				if(in == 3) begin
					state<=4310;
					out<=211;
				end
				if(in == 4) begin
					state<=412;
					out<=212;
				end
			end
			6289: begin
				if(in == 0) begin
					state<=6300;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=2411;
					out<=215;
				end
				if(in == 3) begin
					state<=4311;
					out<=216;
				end
				if(in == 4) begin
					state<=413;
					out<=217;
				end
			end
			6290: begin
				if(in == 0) begin
					state<=6301;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=2412;
					out<=220;
				end
				if(in == 3) begin
					state<=4312;
					out<=221;
				end
				if(in == 4) begin
					state<=414;
					out<=222;
				end
			end
			6291: begin
				if(in == 0) begin
					state<=6292;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=2403;
					out<=225;
				end
				if(in == 3) begin
					state<=4303;
					out<=226;
				end
				if(in == 4) begin
					state<=405;
					out<=227;
				end
			end
			6292: begin
				if(in == 0) begin
					state<=6303;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=2414;
					out<=230;
				end
				if(in == 3) begin
					state<=4314;
					out<=231;
				end
				if(in == 4) begin
					state<=416;
					out<=232;
				end
			end
			6293: begin
				if(in == 0) begin
					state<=6304;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=2415;
					out<=235;
				end
				if(in == 3) begin
					state<=4315;
					out<=236;
				end
				if(in == 4) begin
					state<=417;
					out<=237;
				end
			end
			6294: begin
				if(in == 0) begin
					state<=6305;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=2416;
					out<=240;
				end
				if(in == 3) begin
					state<=4316;
					out<=241;
				end
				if(in == 4) begin
					state<=418;
					out<=242;
				end
			end
			6295: begin
				if(in == 0) begin
					state<=6306;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=2417;
					out<=245;
				end
				if(in == 3) begin
					state<=4317;
					out<=246;
				end
				if(in == 4) begin
					state<=419;
					out<=247;
				end
			end
			6296: begin
				if(in == 0) begin
					state<=6307;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=2418;
					out<=250;
				end
				if(in == 3) begin
					state<=4318;
					out<=251;
				end
				if(in == 4) begin
					state<=420;
					out<=252;
				end
			end
			6297: begin
				if(in == 0) begin
					state<=6308;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=2419;
					out<=255;
				end
				if(in == 3) begin
					state<=4319;
					out<=0;
				end
				if(in == 4) begin
					state<=421;
					out<=1;
				end
			end
			6298: begin
				if(in == 0) begin
					state<=6309;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=2420;
					out<=4;
				end
				if(in == 3) begin
					state<=4320;
					out<=5;
				end
				if(in == 4) begin
					state<=422;
					out<=6;
				end
			end
			6299: begin
				if(in == 0) begin
					state<=6310;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=2421;
					out<=9;
				end
				if(in == 3) begin
					state<=4321;
					out<=10;
				end
				if(in == 4) begin
					state<=423;
					out<=11;
				end
			end
			6300: begin
				if(in == 0) begin
					state<=6311;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=2422;
					out<=14;
				end
				if(in == 3) begin
					state<=4322;
					out<=15;
				end
				if(in == 4) begin
					state<=424;
					out<=16;
				end
			end
			6301: begin
				if(in == 0) begin
					state<=6302;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=2413;
					out<=19;
				end
				if(in == 3) begin
					state<=4313;
					out<=20;
				end
				if(in == 4) begin
					state<=415;
					out<=21;
				end
			end
			6302: begin
				if(in == 0) begin
					state<=6313;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=2424;
					out<=24;
				end
				if(in == 3) begin
					state<=4324;
					out<=25;
				end
				if(in == 4) begin
					state<=426;
					out<=26;
				end
			end
			6303: begin
				if(in == 0) begin
					state<=6314;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=2425;
					out<=29;
				end
				if(in == 3) begin
					state<=4325;
					out<=30;
				end
				if(in == 4) begin
					state<=427;
					out<=31;
				end
			end
			6304: begin
				if(in == 0) begin
					state<=6315;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=2426;
					out<=34;
				end
				if(in == 3) begin
					state<=4326;
					out<=35;
				end
				if(in == 4) begin
					state<=428;
					out<=36;
				end
			end
			6305: begin
				if(in == 0) begin
					state<=6316;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=2427;
					out<=39;
				end
				if(in == 3) begin
					state<=4327;
					out<=40;
				end
				if(in == 4) begin
					state<=429;
					out<=41;
				end
			end
			6306: begin
				if(in == 0) begin
					state<=6317;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=2428;
					out<=44;
				end
				if(in == 3) begin
					state<=4328;
					out<=45;
				end
				if(in == 4) begin
					state<=430;
					out<=46;
				end
			end
			6307: begin
				if(in == 0) begin
					state<=6318;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=2429;
					out<=49;
				end
				if(in == 3) begin
					state<=4329;
					out<=50;
				end
				if(in == 4) begin
					state<=431;
					out<=51;
				end
			end
			6308: begin
				if(in == 0) begin
					state<=6319;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=2430;
					out<=54;
				end
				if(in == 3) begin
					state<=4330;
					out<=55;
				end
				if(in == 4) begin
					state<=432;
					out<=56;
				end
			end
			6309: begin
				if(in == 0) begin
					state<=6320;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=2431;
					out<=59;
				end
				if(in == 3) begin
					state<=4331;
					out<=60;
				end
				if(in == 4) begin
					state<=433;
					out<=61;
				end
			end
			6310: begin
				if(in == 0) begin
					state<=6321;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=2432;
					out<=64;
				end
				if(in == 3) begin
					state<=4332;
					out<=65;
				end
				if(in == 4) begin
					state<=434;
					out<=66;
				end
			end
			6311: begin
				if(in == 0) begin
					state<=6312;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=2423;
					out<=69;
				end
				if(in == 3) begin
					state<=4323;
					out<=70;
				end
				if(in == 4) begin
					state<=425;
					out<=71;
				end
			end
			6312: begin
				if(in == 0) begin
					state<=6323;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=2434;
					out<=74;
				end
				if(in == 3) begin
					state<=4334;
					out<=75;
				end
				if(in == 4) begin
					state<=436;
					out<=76;
				end
			end
			6313: begin
				if(in == 0) begin
					state<=6324;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=2435;
					out<=79;
				end
				if(in == 3) begin
					state<=4335;
					out<=80;
				end
				if(in == 4) begin
					state<=437;
					out<=81;
				end
			end
			6314: begin
				if(in == 0) begin
					state<=6325;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=2436;
					out<=84;
				end
				if(in == 3) begin
					state<=4336;
					out<=85;
				end
				if(in == 4) begin
					state<=438;
					out<=86;
				end
			end
			6315: begin
				if(in == 0) begin
					state<=6326;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=2437;
					out<=89;
				end
				if(in == 3) begin
					state<=4337;
					out<=90;
				end
				if(in == 4) begin
					state<=439;
					out<=91;
				end
			end
			6316: begin
				if(in == 0) begin
					state<=6327;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=2438;
					out<=94;
				end
				if(in == 3) begin
					state<=4338;
					out<=95;
				end
				if(in == 4) begin
					state<=440;
					out<=96;
				end
			end
			6317: begin
				if(in == 0) begin
					state<=6328;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=2439;
					out<=99;
				end
				if(in == 3) begin
					state<=4339;
					out<=100;
				end
				if(in == 4) begin
					state<=441;
					out<=101;
				end
			end
			6318: begin
				if(in == 0) begin
					state<=6329;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=2440;
					out<=104;
				end
				if(in == 3) begin
					state<=4340;
					out<=105;
				end
				if(in == 4) begin
					state<=442;
					out<=106;
				end
			end
			6319: begin
				if(in == 0) begin
					state<=6330;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=2441;
					out<=109;
				end
				if(in == 3) begin
					state<=4341;
					out<=110;
				end
				if(in == 4) begin
					state<=443;
					out<=111;
				end
			end
			6320: begin
				if(in == 0) begin
					state<=6331;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=2442;
					out<=114;
				end
				if(in == 3) begin
					state<=4342;
					out<=115;
				end
				if(in == 4) begin
					state<=444;
					out<=116;
				end
			end
			6321: begin
				if(in == 0) begin
					state<=6322;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=2433;
					out<=119;
				end
				if(in == 3) begin
					state<=4333;
					out<=120;
				end
				if(in == 4) begin
					state<=435;
					out<=121;
				end
			end
			6322: begin
				if(in == 0) begin
					state<=6333;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=2444;
					out<=124;
				end
				if(in == 3) begin
					state<=4344;
					out<=125;
				end
				if(in == 4) begin
					state<=446;
					out<=126;
				end
			end
			6323: begin
				if(in == 0) begin
					state<=6334;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=2445;
					out<=129;
				end
				if(in == 3) begin
					state<=4345;
					out<=130;
				end
				if(in == 4) begin
					state<=447;
					out<=131;
				end
			end
			6324: begin
				if(in == 0) begin
					state<=6335;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=2446;
					out<=134;
				end
				if(in == 3) begin
					state<=4346;
					out<=135;
				end
				if(in == 4) begin
					state<=448;
					out<=136;
				end
			end
			6325: begin
				if(in == 0) begin
					state<=6336;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=2447;
					out<=139;
				end
				if(in == 3) begin
					state<=4347;
					out<=140;
				end
				if(in == 4) begin
					state<=449;
					out<=141;
				end
			end
			6326: begin
				if(in == 0) begin
					state<=6337;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=2448;
					out<=144;
				end
				if(in == 3) begin
					state<=4348;
					out<=145;
				end
				if(in == 4) begin
					state<=450;
					out<=146;
				end
			end
			6327: begin
				if(in == 0) begin
					state<=6338;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=2449;
					out<=149;
				end
				if(in == 3) begin
					state<=4349;
					out<=150;
				end
				if(in == 4) begin
					state<=451;
					out<=151;
				end
			end
			6328: begin
				if(in == 0) begin
					state<=6339;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=2450;
					out<=154;
				end
				if(in == 3) begin
					state<=4350;
					out<=155;
				end
				if(in == 4) begin
					state<=452;
					out<=156;
				end
			end
			6329: begin
				if(in == 0) begin
					state<=6340;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=2451;
					out<=159;
				end
				if(in == 3) begin
					state<=4351;
					out<=160;
				end
				if(in == 4) begin
					state<=453;
					out<=161;
				end
			end
			6330: begin
				if(in == 0) begin
					state<=6341;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=2452;
					out<=164;
				end
				if(in == 3) begin
					state<=4352;
					out<=165;
				end
				if(in == 4) begin
					state<=454;
					out<=166;
				end
			end
			6331: begin
				if(in == 0) begin
					state<=6332;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=2443;
					out<=169;
				end
				if(in == 3) begin
					state<=4343;
					out<=170;
				end
				if(in == 4) begin
					state<=445;
					out<=171;
				end
			end
			6332: begin
				if(in == 0) begin
					state<=6343;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=2454;
					out<=174;
				end
				if(in == 3) begin
					state<=4354;
					out<=175;
				end
				if(in == 4) begin
					state<=456;
					out<=176;
				end
			end
			6333: begin
				if(in == 0) begin
					state<=6344;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=2455;
					out<=179;
				end
				if(in == 3) begin
					state<=4355;
					out<=180;
				end
				if(in == 4) begin
					state<=457;
					out<=181;
				end
			end
			6334: begin
				if(in == 0) begin
					state<=6345;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=2456;
					out<=184;
				end
				if(in == 3) begin
					state<=4356;
					out<=185;
				end
				if(in == 4) begin
					state<=458;
					out<=186;
				end
			end
			6335: begin
				if(in == 0) begin
					state<=6346;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=2457;
					out<=189;
				end
				if(in == 3) begin
					state<=4357;
					out<=190;
				end
				if(in == 4) begin
					state<=459;
					out<=191;
				end
			end
			6336: begin
				if(in == 0) begin
					state<=6347;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=2458;
					out<=194;
				end
				if(in == 3) begin
					state<=4358;
					out<=195;
				end
				if(in == 4) begin
					state<=460;
					out<=196;
				end
			end
			6337: begin
				if(in == 0) begin
					state<=6348;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=2459;
					out<=199;
				end
				if(in == 3) begin
					state<=4359;
					out<=200;
				end
				if(in == 4) begin
					state<=461;
					out<=201;
				end
			end
			6338: begin
				if(in == 0) begin
					state<=6349;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=2460;
					out<=204;
				end
				if(in == 3) begin
					state<=4360;
					out<=205;
				end
				if(in == 4) begin
					state<=462;
					out<=206;
				end
			end
			6339: begin
				if(in == 0) begin
					state<=6350;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=2461;
					out<=209;
				end
				if(in == 3) begin
					state<=4361;
					out<=210;
				end
				if(in == 4) begin
					state<=463;
					out<=211;
				end
			end
			6340: begin
				if(in == 0) begin
					state<=6351;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=2462;
					out<=214;
				end
				if(in == 3) begin
					state<=4362;
					out<=215;
				end
				if(in == 4) begin
					state<=464;
					out<=216;
				end
			end
			6341: begin
				if(in == 0) begin
					state<=6342;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=2453;
					out<=219;
				end
				if(in == 3) begin
					state<=4353;
					out<=220;
				end
				if(in == 4) begin
					state<=455;
					out<=221;
				end
			end
			6342: begin
				if(in == 0) begin
					state<=7306;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=3417;
					out<=224;
				end
				if(in == 3) begin
					state<=5374;
					out<=225;
				end
				if(in == 4) begin
					state<=1485;
					out<=226;
				end
			end
			6343: begin
				if(in == 0) begin
					state<=7307;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=3418;
					out<=229;
				end
				if(in == 3) begin
					state<=5375;
					out<=230;
				end
				if(in == 4) begin
					state<=1486;
					out<=231;
				end
			end
			6344: begin
				if(in == 0) begin
					state<=7308;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=3419;
					out<=234;
				end
				if(in == 3) begin
					state<=5376;
					out<=235;
				end
				if(in == 4) begin
					state<=1487;
					out<=236;
				end
			end
			6345: begin
				if(in == 0) begin
					state<=7309;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=3420;
					out<=239;
				end
				if(in == 3) begin
					state<=5377;
					out<=240;
				end
				if(in == 4) begin
					state<=1488;
					out<=241;
				end
			end
			6346: begin
				if(in == 0) begin
					state<=7310;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=3421;
					out<=244;
				end
				if(in == 3) begin
					state<=5378;
					out<=245;
				end
				if(in == 4) begin
					state<=1489;
					out<=246;
				end
			end
			6347: begin
				if(in == 0) begin
					state<=7311;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=3422;
					out<=249;
				end
				if(in == 3) begin
					state<=5379;
					out<=250;
				end
				if(in == 4) begin
					state<=1490;
					out<=251;
				end
			end
			6348: begin
				if(in == 0) begin
					state<=7312;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=3423;
					out<=254;
				end
				if(in == 3) begin
					state<=5380;
					out<=255;
				end
				if(in == 4) begin
					state<=1491;
					out<=0;
				end
			end
			6349: begin
				if(in == 0) begin
					state<=7313;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=3424;
					out<=3;
				end
				if(in == 3) begin
					state<=5381;
					out<=4;
				end
				if(in == 4) begin
					state<=1492;
					out<=5;
				end
			end
			6350: begin
				if(in == 0) begin
					state<=7314;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=3425;
					out<=8;
				end
				if(in == 3) begin
					state<=5382;
					out<=9;
				end
				if(in == 4) begin
					state<=1493;
					out<=10;
				end
			end
			6351: begin
				if(in == 0) begin
					state<=7305;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=3416;
					out<=13;
				end
				if(in == 3) begin
					state<=5373;
					out<=14;
				end
				if(in == 4) begin
					state<=1484;
					out<=15;
				end
			end
			6352: begin
				if(in == 0) begin
					state<=6363;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=2474;
					out<=18;
				end
				if(in == 3) begin
					state<=4374;
					out<=19;
				end
				if(in == 4) begin
					state<=476;
					out<=20;
				end
			end
			6353: begin
				if(in == 0) begin
					state<=6364;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=2475;
					out<=23;
				end
				if(in == 3) begin
					state<=4375;
					out<=24;
				end
				if(in == 4) begin
					state<=477;
					out<=25;
				end
			end
			6354: begin
				if(in == 0) begin
					state<=6365;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=2476;
					out<=28;
				end
				if(in == 3) begin
					state<=4376;
					out<=29;
				end
				if(in == 4) begin
					state<=478;
					out<=30;
				end
			end
			6355: begin
				if(in == 0) begin
					state<=6366;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=2477;
					out<=33;
				end
				if(in == 3) begin
					state<=4377;
					out<=34;
				end
				if(in == 4) begin
					state<=479;
					out<=35;
				end
			end
			6356: begin
				if(in == 0) begin
					state<=6367;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=2478;
					out<=38;
				end
				if(in == 3) begin
					state<=4378;
					out<=39;
				end
				if(in == 4) begin
					state<=480;
					out<=40;
				end
			end
			6357: begin
				if(in == 0) begin
					state<=6368;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=2479;
					out<=43;
				end
				if(in == 3) begin
					state<=4379;
					out<=44;
				end
				if(in == 4) begin
					state<=481;
					out<=45;
				end
			end
			6358: begin
				if(in == 0) begin
					state<=6369;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=2480;
					out<=48;
				end
				if(in == 3) begin
					state<=4380;
					out<=49;
				end
				if(in == 4) begin
					state<=482;
					out<=50;
				end
			end
			6359: begin
				if(in == 0) begin
					state<=6370;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=2481;
					out<=53;
				end
				if(in == 3) begin
					state<=4381;
					out<=54;
				end
				if(in == 4) begin
					state<=483;
					out<=55;
				end
			end
			6360: begin
				if(in == 0) begin
					state<=6361;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=2472;
					out<=58;
				end
				if(in == 3) begin
					state<=4372;
					out<=59;
				end
				if(in == 4) begin
					state<=474;
					out<=60;
				end
			end
			6361: begin
				if(in == 0) begin
					state<=6372;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=2483;
					out<=63;
				end
				if(in == 3) begin
					state<=4383;
					out<=64;
				end
				if(in == 4) begin
					state<=485;
					out<=65;
				end
			end
			6362: begin
				if(in == 0) begin
					state<=6373;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=2484;
					out<=68;
				end
				if(in == 3) begin
					state<=4384;
					out<=69;
				end
				if(in == 4) begin
					state<=486;
					out<=70;
				end
			end
			6363: begin
				if(in == 0) begin
					state<=6374;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=2485;
					out<=73;
				end
				if(in == 3) begin
					state<=4385;
					out<=74;
				end
				if(in == 4) begin
					state<=487;
					out<=75;
				end
			end
			6364: begin
				if(in == 0) begin
					state<=6375;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=2486;
					out<=78;
				end
				if(in == 3) begin
					state<=4386;
					out<=79;
				end
				if(in == 4) begin
					state<=488;
					out<=80;
				end
			end
			6365: begin
				if(in == 0) begin
					state<=6376;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=2487;
					out<=83;
				end
				if(in == 3) begin
					state<=4387;
					out<=84;
				end
				if(in == 4) begin
					state<=489;
					out<=85;
				end
			end
			6366: begin
				if(in == 0) begin
					state<=6377;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=2488;
					out<=88;
				end
				if(in == 3) begin
					state<=4388;
					out<=89;
				end
				if(in == 4) begin
					state<=490;
					out<=90;
				end
			end
			6367: begin
				if(in == 0) begin
					state<=6378;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=2489;
					out<=93;
				end
				if(in == 3) begin
					state<=4389;
					out<=94;
				end
				if(in == 4) begin
					state<=491;
					out<=95;
				end
			end
			6368: begin
				if(in == 0) begin
					state<=6379;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=2490;
					out<=98;
				end
				if(in == 3) begin
					state<=4390;
					out<=99;
				end
				if(in == 4) begin
					state<=492;
					out<=100;
				end
			end
			6369: begin
				if(in == 0) begin
					state<=6380;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=2491;
					out<=103;
				end
				if(in == 3) begin
					state<=4391;
					out<=104;
				end
				if(in == 4) begin
					state<=493;
					out<=105;
				end
			end
			6370: begin
				if(in == 0) begin
					state<=6371;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=2482;
					out<=108;
				end
				if(in == 3) begin
					state<=4382;
					out<=109;
				end
				if(in == 4) begin
					state<=484;
					out<=110;
				end
			end
			6371: begin
				if(in == 0) begin
					state<=6382;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=2493;
					out<=113;
				end
				if(in == 3) begin
					state<=4393;
					out<=114;
				end
				if(in == 4) begin
					state<=495;
					out<=115;
				end
			end
			6372: begin
				if(in == 0) begin
					state<=6383;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=2494;
					out<=118;
				end
				if(in == 3) begin
					state<=4394;
					out<=119;
				end
				if(in == 4) begin
					state<=496;
					out<=120;
				end
			end
			6373: begin
				if(in == 0) begin
					state<=6384;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=2495;
					out<=123;
				end
				if(in == 3) begin
					state<=4395;
					out<=124;
				end
				if(in == 4) begin
					state<=497;
					out<=125;
				end
			end
			6374: begin
				if(in == 0) begin
					state<=6385;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=2496;
					out<=128;
				end
				if(in == 3) begin
					state<=4396;
					out<=129;
				end
				if(in == 4) begin
					state<=498;
					out<=130;
				end
			end
			6375: begin
				if(in == 0) begin
					state<=6386;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=2497;
					out<=133;
				end
				if(in == 3) begin
					state<=4397;
					out<=134;
				end
				if(in == 4) begin
					state<=499;
					out<=135;
				end
			end
			6376: begin
				if(in == 0) begin
					state<=6387;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=2498;
					out<=138;
				end
				if(in == 3) begin
					state<=4398;
					out<=139;
				end
				if(in == 4) begin
					state<=500;
					out<=140;
				end
			end
			6377: begin
				if(in == 0) begin
					state<=6388;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=2499;
					out<=143;
				end
				if(in == 3) begin
					state<=4399;
					out<=144;
				end
				if(in == 4) begin
					state<=501;
					out<=145;
				end
			end
			6378: begin
				if(in == 0) begin
					state<=6389;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=2500;
					out<=148;
				end
				if(in == 3) begin
					state<=4400;
					out<=149;
				end
				if(in == 4) begin
					state<=502;
					out<=150;
				end
			end
			6379: begin
				if(in == 0) begin
					state<=6390;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=2501;
					out<=153;
				end
				if(in == 3) begin
					state<=4401;
					out<=154;
				end
				if(in == 4) begin
					state<=503;
					out<=155;
				end
			end
			6380: begin
				if(in == 0) begin
					state<=6381;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=2492;
					out<=158;
				end
				if(in == 3) begin
					state<=4392;
					out<=159;
				end
				if(in == 4) begin
					state<=494;
					out<=160;
				end
			end
			6381: begin
				if(in == 0) begin
					state<=6392;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=2503;
					out<=163;
				end
				if(in == 3) begin
					state<=4403;
					out<=164;
				end
				if(in == 4) begin
					state<=505;
					out<=165;
				end
			end
			6382: begin
				if(in == 0) begin
					state<=6393;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=2504;
					out<=168;
				end
				if(in == 3) begin
					state<=4404;
					out<=169;
				end
				if(in == 4) begin
					state<=506;
					out<=170;
				end
			end
			6383: begin
				if(in == 0) begin
					state<=6394;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=2505;
					out<=173;
				end
				if(in == 3) begin
					state<=4405;
					out<=174;
				end
				if(in == 4) begin
					state<=507;
					out<=175;
				end
			end
			6384: begin
				if(in == 0) begin
					state<=6395;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=2506;
					out<=178;
				end
				if(in == 3) begin
					state<=4406;
					out<=179;
				end
				if(in == 4) begin
					state<=508;
					out<=180;
				end
			end
			6385: begin
				if(in == 0) begin
					state<=6396;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=2507;
					out<=183;
				end
				if(in == 3) begin
					state<=4407;
					out<=184;
				end
				if(in == 4) begin
					state<=509;
					out<=185;
				end
			end
			6386: begin
				if(in == 0) begin
					state<=6397;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=2508;
					out<=188;
				end
				if(in == 3) begin
					state<=4408;
					out<=189;
				end
				if(in == 4) begin
					state<=510;
					out<=190;
				end
			end
			6387: begin
				if(in == 0) begin
					state<=6398;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=2509;
					out<=193;
				end
				if(in == 3) begin
					state<=4409;
					out<=194;
				end
				if(in == 4) begin
					state<=511;
					out<=195;
				end
			end
			6388: begin
				if(in == 0) begin
					state<=6399;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=2510;
					out<=198;
				end
				if(in == 3) begin
					state<=4410;
					out<=199;
				end
				if(in == 4) begin
					state<=512;
					out<=200;
				end
			end
			6389: begin
				if(in == 0) begin
					state<=6400;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=2511;
					out<=203;
				end
				if(in == 3) begin
					state<=4411;
					out<=204;
				end
				if(in == 4) begin
					state<=513;
					out<=205;
				end
			end
			6390: begin
				if(in == 0) begin
					state<=6391;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=2502;
					out<=208;
				end
				if(in == 3) begin
					state<=4402;
					out<=209;
				end
				if(in == 4) begin
					state<=504;
					out<=210;
				end
			end
			6391: begin
				if(in == 0) begin
					state<=6402;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=2513;
					out<=213;
				end
				if(in == 3) begin
					state<=4413;
					out<=214;
				end
				if(in == 4) begin
					state<=515;
					out<=215;
				end
			end
			6392: begin
				if(in == 0) begin
					state<=6403;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=2514;
					out<=218;
				end
				if(in == 3) begin
					state<=4414;
					out<=219;
				end
				if(in == 4) begin
					state<=516;
					out<=220;
				end
			end
			6393: begin
				if(in == 0) begin
					state<=6404;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=2515;
					out<=223;
				end
				if(in == 3) begin
					state<=4415;
					out<=224;
				end
				if(in == 4) begin
					state<=517;
					out<=225;
				end
			end
			6394: begin
				if(in == 0) begin
					state<=6405;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=2516;
					out<=228;
				end
				if(in == 3) begin
					state<=4416;
					out<=229;
				end
				if(in == 4) begin
					state<=518;
					out<=230;
				end
			end
			6395: begin
				if(in == 0) begin
					state<=6406;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=2517;
					out<=233;
				end
				if(in == 3) begin
					state<=4417;
					out<=234;
				end
				if(in == 4) begin
					state<=519;
					out<=235;
				end
			end
			6396: begin
				if(in == 0) begin
					state<=6407;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=2518;
					out<=238;
				end
				if(in == 3) begin
					state<=4418;
					out<=239;
				end
				if(in == 4) begin
					state<=520;
					out<=240;
				end
			end
			6397: begin
				if(in == 0) begin
					state<=6408;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=2519;
					out<=243;
				end
				if(in == 3) begin
					state<=4419;
					out<=244;
				end
				if(in == 4) begin
					state<=521;
					out<=245;
				end
			end
			6398: begin
				if(in == 0) begin
					state<=6409;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=2520;
					out<=248;
				end
				if(in == 3) begin
					state<=4420;
					out<=249;
				end
				if(in == 4) begin
					state<=522;
					out<=250;
				end
			end
			6399: begin
				if(in == 0) begin
					state<=6410;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=2521;
					out<=253;
				end
				if(in == 3) begin
					state<=4421;
					out<=254;
				end
				if(in == 4) begin
					state<=523;
					out<=255;
				end
			end
			6400: begin
				if(in == 0) begin
					state<=6401;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=2512;
					out<=2;
				end
				if(in == 3) begin
					state<=4412;
					out<=3;
				end
				if(in == 4) begin
					state<=514;
					out<=4;
				end
			end
			6401: begin
				if(in == 0) begin
					state<=6412;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=2523;
					out<=7;
				end
				if(in == 3) begin
					state<=4423;
					out<=8;
				end
				if(in == 4) begin
					state<=525;
					out<=9;
				end
			end
			6402: begin
				if(in == 0) begin
					state<=6413;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=2524;
					out<=12;
				end
				if(in == 3) begin
					state<=4424;
					out<=13;
				end
				if(in == 4) begin
					state<=526;
					out<=14;
				end
			end
			6403: begin
				if(in == 0) begin
					state<=6414;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=2525;
					out<=17;
				end
				if(in == 3) begin
					state<=4425;
					out<=18;
				end
				if(in == 4) begin
					state<=527;
					out<=19;
				end
			end
			6404: begin
				if(in == 0) begin
					state<=6415;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=2526;
					out<=22;
				end
				if(in == 3) begin
					state<=4426;
					out<=23;
				end
				if(in == 4) begin
					state<=528;
					out<=24;
				end
			end
			6405: begin
				if(in == 0) begin
					state<=6416;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=2527;
					out<=27;
				end
				if(in == 3) begin
					state<=4427;
					out<=28;
				end
				if(in == 4) begin
					state<=529;
					out<=29;
				end
			end
			6406: begin
				if(in == 0) begin
					state<=6417;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=2528;
					out<=32;
				end
				if(in == 3) begin
					state<=4428;
					out<=33;
				end
				if(in == 4) begin
					state<=530;
					out<=34;
				end
			end
			6407: begin
				if(in == 0) begin
					state<=6418;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=2529;
					out<=37;
				end
				if(in == 3) begin
					state<=4429;
					out<=38;
				end
				if(in == 4) begin
					state<=531;
					out<=39;
				end
			end
			6408: begin
				if(in == 0) begin
					state<=6419;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=2530;
					out<=42;
				end
				if(in == 3) begin
					state<=4430;
					out<=43;
				end
				if(in == 4) begin
					state<=532;
					out<=44;
				end
			end
			6409: begin
				if(in == 0) begin
					state<=6420;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=2531;
					out<=47;
				end
				if(in == 3) begin
					state<=4431;
					out<=48;
				end
				if(in == 4) begin
					state<=533;
					out<=49;
				end
			end
			6410: begin
				if(in == 0) begin
					state<=6411;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=2522;
					out<=52;
				end
				if(in == 3) begin
					state<=4422;
					out<=53;
				end
				if(in == 4) begin
					state<=524;
					out<=54;
				end
			end
			6411: begin
				if(in == 0) begin
					state<=7337;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=3448;
					out<=57;
				end
				if(in == 3) begin
					state<=5405;
					out<=58;
				end
				if(in == 4) begin
					state<=1516;
					out<=59;
				end
			end
			6412: begin
				if(in == 0) begin
					state<=7338;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=3449;
					out<=62;
				end
				if(in == 3) begin
					state<=5406;
					out<=63;
				end
				if(in == 4) begin
					state<=1517;
					out<=64;
				end
			end
			6413: begin
				if(in == 0) begin
					state<=7339;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=3450;
					out<=67;
				end
				if(in == 3) begin
					state<=5407;
					out<=68;
				end
				if(in == 4) begin
					state<=1518;
					out<=69;
				end
			end
			6414: begin
				if(in == 0) begin
					state<=7340;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=3451;
					out<=72;
				end
				if(in == 3) begin
					state<=5408;
					out<=73;
				end
				if(in == 4) begin
					state<=1519;
					out<=74;
				end
			end
			6415: begin
				if(in == 0) begin
					state<=7341;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=3452;
					out<=77;
				end
				if(in == 3) begin
					state<=5409;
					out<=78;
				end
				if(in == 4) begin
					state<=1520;
					out<=79;
				end
			end
			6416: begin
				if(in == 0) begin
					state<=7342;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=3453;
					out<=82;
				end
				if(in == 3) begin
					state<=5410;
					out<=83;
				end
				if(in == 4) begin
					state<=1521;
					out<=84;
				end
			end
			6417: begin
				if(in == 0) begin
					state<=7343;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=3454;
					out<=87;
				end
				if(in == 3) begin
					state<=5411;
					out<=88;
				end
				if(in == 4) begin
					state<=1522;
					out<=89;
				end
			end
			6418: begin
				if(in == 0) begin
					state<=7344;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=3455;
					out<=92;
				end
				if(in == 3) begin
					state<=5412;
					out<=93;
				end
				if(in == 4) begin
					state<=1523;
					out<=94;
				end
			end
			6419: begin
				if(in == 0) begin
					state<=7345;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=3456;
					out<=97;
				end
				if(in == 3) begin
					state<=5413;
					out<=98;
				end
				if(in == 4) begin
					state<=1524;
					out<=99;
				end
			end
			6420: begin
				if(in == 0) begin
					state<=7336;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=3447;
					out<=102;
				end
				if(in == 3) begin
					state<=5404;
					out<=103;
				end
				if(in == 4) begin
					state<=1515;
					out<=104;
				end
			end
			6421: begin
				if(in == 0) begin
					state<=6432;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=2543;
					out<=107;
				end
				if(in == 3) begin
					state<=4443;
					out<=108;
				end
				if(in == 4) begin
					state<=545;
					out<=109;
				end
			end
			6422: begin
				if(in == 0) begin
					state<=6433;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=2544;
					out<=112;
				end
				if(in == 3) begin
					state<=4444;
					out<=113;
				end
				if(in == 4) begin
					state<=546;
					out<=114;
				end
			end
			6423: begin
				if(in == 0) begin
					state<=6434;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=2545;
					out<=117;
				end
				if(in == 3) begin
					state<=4445;
					out<=118;
				end
				if(in == 4) begin
					state<=547;
					out<=119;
				end
			end
			6424: begin
				if(in == 0) begin
					state<=6435;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=2546;
					out<=122;
				end
				if(in == 3) begin
					state<=4446;
					out<=123;
				end
				if(in == 4) begin
					state<=548;
					out<=124;
				end
			end
			6425: begin
				if(in == 0) begin
					state<=6436;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=2547;
					out<=127;
				end
				if(in == 3) begin
					state<=4447;
					out<=128;
				end
				if(in == 4) begin
					state<=549;
					out<=129;
				end
			end
			6426: begin
				if(in == 0) begin
					state<=6437;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=2548;
					out<=132;
				end
				if(in == 3) begin
					state<=4448;
					out<=133;
				end
				if(in == 4) begin
					state<=550;
					out<=134;
				end
			end
			6427: begin
				if(in == 0) begin
					state<=6438;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=2549;
					out<=137;
				end
				if(in == 3) begin
					state<=4449;
					out<=138;
				end
				if(in == 4) begin
					state<=551;
					out<=139;
				end
			end
			6428: begin
				if(in == 0) begin
					state<=6439;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=2550;
					out<=142;
				end
				if(in == 3) begin
					state<=4450;
					out<=143;
				end
				if(in == 4) begin
					state<=552;
					out<=144;
				end
			end
			6429: begin
				if(in == 0) begin
					state<=6430;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=2541;
					out<=147;
				end
				if(in == 3) begin
					state<=4441;
					out<=148;
				end
				if(in == 4) begin
					state<=543;
					out<=149;
				end
			end
			6430: begin
				if(in == 0) begin
					state<=6441;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=2552;
					out<=152;
				end
				if(in == 3) begin
					state<=4452;
					out<=153;
				end
				if(in == 4) begin
					state<=554;
					out<=154;
				end
			end
			6431: begin
				if(in == 0) begin
					state<=6442;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=2553;
					out<=157;
				end
				if(in == 3) begin
					state<=4453;
					out<=158;
				end
				if(in == 4) begin
					state<=555;
					out<=159;
				end
			end
			6432: begin
				if(in == 0) begin
					state<=6443;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=2554;
					out<=162;
				end
				if(in == 3) begin
					state<=4454;
					out<=163;
				end
				if(in == 4) begin
					state<=556;
					out<=164;
				end
			end
			6433: begin
				if(in == 0) begin
					state<=6444;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=2555;
					out<=167;
				end
				if(in == 3) begin
					state<=4455;
					out<=168;
				end
				if(in == 4) begin
					state<=557;
					out<=169;
				end
			end
			6434: begin
				if(in == 0) begin
					state<=6445;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=2556;
					out<=172;
				end
				if(in == 3) begin
					state<=4456;
					out<=173;
				end
				if(in == 4) begin
					state<=558;
					out<=174;
				end
			end
			6435: begin
				if(in == 0) begin
					state<=6446;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=2557;
					out<=177;
				end
				if(in == 3) begin
					state<=4457;
					out<=178;
				end
				if(in == 4) begin
					state<=559;
					out<=179;
				end
			end
			6436: begin
				if(in == 0) begin
					state<=6447;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=2558;
					out<=182;
				end
				if(in == 3) begin
					state<=4458;
					out<=183;
				end
				if(in == 4) begin
					state<=560;
					out<=184;
				end
			end
			6437: begin
				if(in == 0) begin
					state<=6448;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=2559;
					out<=187;
				end
				if(in == 3) begin
					state<=4459;
					out<=188;
				end
				if(in == 4) begin
					state<=561;
					out<=189;
				end
			end
			6438: begin
				if(in == 0) begin
					state<=6449;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=2560;
					out<=192;
				end
				if(in == 3) begin
					state<=4460;
					out<=193;
				end
				if(in == 4) begin
					state<=562;
					out<=194;
				end
			end
			6439: begin
				if(in == 0) begin
					state<=6440;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=2551;
					out<=197;
				end
				if(in == 3) begin
					state<=4451;
					out<=198;
				end
				if(in == 4) begin
					state<=553;
					out<=199;
				end
			end
			6440: begin
				if(in == 0) begin
					state<=6451;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=2562;
					out<=202;
				end
				if(in == 3) begin
					state<=4462;
					out<=203;
				end
				if(in == 4) begin
					state<=564;
					out<=204;
				end
			end
			6441: begin
				if(in == 0) begin
					state<=6452;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=2563;
					out<=207;
				end
				if(in == 3) begin
					state<=4463;
					out<=208;
				end
				if(in == 4) begin
					state<=565;
					out<=209;
				end
			end
			6442: begin
				if(in == 0) begin
					state<=6453;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=2564;
					out<=212;
				end
				if(in == 3) begin
					state<=4464;
					out<=213;
				end
				if(in == 4) begin
					state<=566;
					out<=214;
				end
			end
			6443: begin
				if(in == 0) begin
					state<=6454;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=2565;
					out<=217;
				end
				if(in == 3) begin
					state<=4465;
					out<=218;
				end
				if(in == 4) begin
					state<=567;
					out<=219;
				end
			end
			6444: begin
				if(in == 0) begin
					state<=6455;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=2566;
					out<=222;
				end
				if(in == 3) begin
					state<=4466;
					out<=223;
				end
				if(in == 4) begin
					state<=568;
					out<=224;
				end
			end
			6445: begin
				if(in == 0) begin
					state<=6456;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=2567;
					out<=227;
				end
				if(in == 3) begin
					state<=4467;
					out<=228;
				end
				if(in == 4) begin
					state<=569;
					out<=229;
				end
			end
			6446: begin
				if(in == 0) begin
					state<=6457;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=2568;
					out<=232;
				end
				if(in == 3) begin
					state<=4468;
					out<=233;
				end
				if(in == 4) begin
					state<=570;
					out<=234;
				end
			end
			6447: begin
				if(in == 0) begin
					state<=6458;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=2569;
					out<=237;
				end
				if(in == 3) begin
					state<=4469;
					out<=238;
				end
				if(in == 4) begin
					state<=571;
					out<=239;
				end
			end
			6448: begin
				if(in == 0) begin
					state<=6459;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=2570;
					out<=242;
				end
				if(in == 3) begin
					state<=4470;
					out<=243;
				end
				if(in == 4) begin
					state<=572;
					out<=244;
				end
			end
			6449: begin
				if(in == 0) begin
					state<=6450;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=2561;
					out<=247;
				end
				if(in == 3) begin
					state<=4461;
					out<=248;
				end
				if(in == 4) begin
					state<=563;
					out<=249;
				end
			end
			6450: begin
				if(in == 0) begin
					state<=6461;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=2572;
					out<=252;
				end
				if(in == 3) begin
					state<=4472;
					out<=253;
				end
				if(in == 4) begin
					state<=574;
					out<=254;
				end
			end
			6451: begin
				if(in == 0) begin
					state<=6462;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=2573;
					out<=1;
				end
				if(in == 3) begin
					state<=4473;
					out<=2;
				end
				if(in == 4) begin
					state<=575;
					out<=3;
				end
			end
			6452: begin
				if(in == 0) begin
					state<=6463;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=2574;
					out<=6;
				end
				if(in == 3) begin
					state<=4474;
					out<=7;
				end
				if(in == 4) begin
					state<=576;
					out<=8;
				end
			end
			6453: begin
				if(in == 0) begin
					state<=6464;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=2575;
					out<=11;
				end
				if(in == 3) begin
					state<=4475;
					out<=12;
				end
				if(in == 4) begin
					state<=577;
					out<=13;
				end
			end
			6454: begin
				if(in == 0) begin
					state<=6465;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=2576;
					out<=16;
				end
				if(in == 3) begin
					state<=4476;
					out<=17;
				end
				if(in == 4) begin
					state<=578;
					out<=18;
				end
			end
			6455: begin
				if(in == 0) begin
					state<=6466;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=2577;
					out<=21;
				end
				if(in == 3) begin
					state<=4477;
					out<=22;
				end
				if(in == 4) begin
					state<=579;
					out<=23;
				end
			end
			6456: begin
				if(in == 0) begin
					state<=6467;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=2578;
					out<=26;
				end
				if(in == 3) begin
					state<=4478;
					out<=27;
				end
				if(in == 4) begin
					state<=580;
					out<=28;
				end
			end
			6457: begin
				if(in == 0) begin
					state<=6468;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=2579;
					out<=31;
				end
				if(in == 3) begin
					state<=4479;
					out<=32;
				end
				if(in == 4) begin
					state<=581;
					out<=33;
				end
			end
			6458: begin
				if(in == 0) begin
					state<=6469;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=2580;
					out<=36;
				end
				if(in == 3) begin
					state<=4480;
					out<=37;
				end
				if(in == 4) begin
					state<=582;
					out<=38;
				end
			end
			6459: begin
				if(in == 0) begin
					state<=6460;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=2571;
					out<=41;
				end
				if(in == 3) begin
					state<=4471;
					out<=42;
				end
				if(in == 4) begin
					state<=573;
					out<=43;
				end
			end
			6460: begin
				if(in == 0) begin
					state<=6471;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=2582;
					out<=46;
				end
				if(in == 3) begin
					state<=4482;
					out<=47;
				end
				if(in == 4) begin
					state<=584;
					out<=48;
				end
			end
			6461: begin
				if(in == 0) begin
					state<=6472;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=2583;
					out<=51;
				end
				if(in == 3) begin
					state<=4483;
					out<=52;
				end
				if(in == 4) begin
					state<=585;
					out<=53;
				end
			end
			6462: begin
				if(in == 0) begin
					state<=6473;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=2584;
					out<=56;
				end
				if(in == 3) begin
					state<=4484;
					out<=57;
				end
				if(in == 4) begin
					state<=586;
					out<=58;
				end
			end
			6463: begin
				if(in == 0) begin
					state<=6474;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=2585;
					out<=61;
				end
				if(in == 3) begin
					state<=4485;
					out<=62;
				end
				if(in == 4) begin
					state<=587;
					out<=63;
				end
			end
			6464: begin
				if(in == 0) begin
					state<=6475;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=2586;
					out<=66;
				end
				if(in == 3) begin
					state<=4486;
					out<=67;
				end
				if(in == 4) begin
					state<=588;
					out<=68;
				end
			end
			6465: begin
				if(in == 0) begin
					state<=6476;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=2587;
					out<=71;
				end
				if(in == 3) begin
					state<=4487;
					out<=72;
				end
				if(in == 4) begin
					state<=589;
					out<=73;
				end
			end
			6466: begin
				if(in == 0) begin
					state<=6477;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=2588;
					out<=76;
				end
				if(in == 3) begin
					state<=4488;
					out<=77;
				end
				if(in == 4) begin
					state<=590;
					out<=78;
				end
			end
			6467: begin
				if(in == 0) begin
					state<=6478;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=2589;
					out<=81;
				end
				if(in == 3) begin
					state<=4489;
					out<=82;
				end
				if(in == 4) begin
					state<=591;
					out<=83;
				end
			end
			6468: begin
				if(in == 0) begin
					state<=6479;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=2590;
					out<=86;
				end
				if(in == 3) begin
					state<=4490;
					out<=87;
				end
				if(in == 4) begin
					state<=592;
					out<=88;
				end
			end
			6469: begin
				if(in == 0) begin
					state<=6470;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=2581;
					out<=91;
				end
				if(in == 3) begin
					state<=4481;
					out<=92;
				end
				if(in == 4) begin
					state<=583;
					out<=93;
				end
			end
			6470: begin
				if(in == 0) begin
					state<=6481;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=2592;
					out<=96;
				end
				if(in == 3) begin
					state<=4492;
					out<=97;
				end
				if(in == 4) begin
					state<=594;
					out<=98;
				end
			end
			6471: begin
				if(in == 0) begin
					state<=6482;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=2593;
					out<=101;
				end
				if(in == 3) begin
					state<=4493;
					out<=102;
				end
				if(in == 4) begin
					state<=595;
					out<=103;
				end
			end
			6472: begin
				if(in == 0) begin
					state<=6483;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=2594;
					out<=106;
				end
				if(in == 3) begin
					state<=4494;
					out<=107;
				end
				if(in == 4) begin
					state<=596;
					out<=108;
				end
			end
			6473: begin
				if(in == 0) begin
					state<=6484;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=2595;
					out<=111;
				end
				if(in == 3) begin
					state<=4495;
					out<=112;
				end
				if(in == 4) begin
					state<=597;
					out<=113;
				end
			end
			6474: begin
				if(in == 0) begin
					state<=6485;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=2596;
					out<=116;
				end
				if(in == 3) begin
					state<=4496;
					out<=117;
				end
				if(in == 4) begin
					state<=598;
					out<=118;
				end
			end
			6475: begin
				if(in == 0) begin
					state<=6486;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=2597;
					out<=121;
				end
				if(in == 3) begin
					state<=4497;
					out<=122;
				end
				if(in == 4) begin
					state<=599;
					out<=123;
				end
			end
			6476: begin
				if(in == 0) begin
					state<=6487;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=2598;
					out<=126;
				end
				if(in == 3) begin
					state<=4498;
					out<=127;
				end
				if(in == 4) begin
					state<=600;
					out<=128;
				end
			end
			6477: begin
				if(in == 0) begin
					state<=6488;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=2599;
					out<=131;
				end
				if(in == 3) begin
					state<=4499;
					out<=132;
				end
				if(in == 4) begin
					state<=601;
					out<=133;
				end
			end
			6478: begin
				if(in == 0) begin
					state<=6489;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=2600;
					out<=136;
				end
				if(in == 3) begin
					state<=4500;
					out<=137;
				end
				if(in == 4) begin
					state<=602;
					out<=138;
				end
			end
			6479: begin
				if(in == 0) begin
					state<=6480;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=2591;
					out<=141;
				end
				if(in == 3) begin
					state<=4491;
					out<=142;
				end
				if(in == 4) begin
					state<=593;
					out<=143;
				end
			end
			6480: begin
				if(in == 0) begin
					state<=7368;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=3479;
					out<=146;
				end
				if(in == 3) begin
					state<=5436;
					out<=147;
				end
				if(in == 4) begin
					state<=1547;
					out<=148;
				end
			end
			6481: begin
				if(in == 0) begin
					state<=7369;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=3480;
					out<=151;
				end
				if(in == 3) begin
					state<=5437;
					out<=152;
				end
				if(in == 4) begin
					state<=1548;
					out<=153;
				end
			end
			6482: begin
				if(in == 0) begin
					state<=7370;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=3481;
					out<=156;
				end
				if(in == 3) begin
					state<=5438;
					out<=157;
				end
				if(in == 4) begin
					state<=1549;
					out<=158;
				end
			end
			6483: begin
				if(in == 0) begin
					state<=7371;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=3482;
					out<=161;
				end
				if(in == 3) begin
					state<=5439;
					out<=162;
				end
				if(in == 4) begin
					state<=1550;
					out<=163;
				end
			end
			6484: begin
				if(in == 0) begin
					state<=7372;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=3483;
					out<=166;
				end
				if(in == 3) begin
					state<=5440;
					out<=167;
				end
				if(in == 4) begin
					state<=1551;
					out<=168;
				end
			end
			6485: begin
				if(in == 0) begin
					state<=7373;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=3484;
					out<=171;
				end
				if(in == 3) begin
					state<=5441;
					out<=172;
				end
				if(in == 4) begin
					state<=1552;
					out<=173;
				end
			end
			6486: begin
				if(in == 0) begin
					state<=7374;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=3485;
					out<=176;
				end
				if(in == 3) begin
					state<=5442;
					out<=177;
				end
				if(in == 4) begin
					state<=1553;
					out<=178;
				end
			end
			6487: begin
				if(in == 0) begin
					state<=7375;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=3486;
					out<=181;
				end
				if(in == 3) begin
					state<=5443;
					out<=182;
				end
				if(in == 4) begin
					state<=1554;
					out<=183;
				end
			end
			6488: begin
				if(in == 0) begin
					state<=7376;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=3487;
					out<=186;
				end
				if(in == 3) begin
					state<=5444;
					out<=187;
				end
				if(in == 4) begin
					state<=1555;
					out<=188;
				end
			end
			6489: begin
				if(in == 0) begin
					state<=7367;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=3478;
					out<=191;
				end
				if(in == 3) begin
					state<=5435;
					out<=192;
				end
				if(in == 4) begin
					state<=1546;
					out<=193;
				end
			end
			6490: begin
				if(in == 0) begin
					state<=6501;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=2612;
					out<=196;
				end
				if(in == 3) begin
					state<=4512;
					out<=197;
				end
				if(in == 4) begin
					state<=614;
					out<=198;
				end
			end
			6491: begin
				if(in == 0) begin
					state<=6502;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=2613;
					out<=201;
				end
				if(in == 3) begin
					state<=4513;
					out<=202;
				end
				if(in == 4) begin
					state<=615;
					out<=203;
				end
			end
			6492: begin
				if(in == 0) begin
					state<=6503;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=2614;
					out<=206;
				end
				if(in == 3) begin
					state<=4514;
					out<=207;
				end
				if(in == 4) begin
					state<=616;
					out<=208;
				end
			end
			6493: begin
				if(in == 0) begin
					state<=6504;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=2615;
					out<=211;
				end
				if(in == 3) begin
					state<=4515;
					out<=212;
				end
				if(in == 4) begin
					state<=617;
					out<=213;
				end
			end
			6494: begin
				if(in == 0) begin
					state<=6505;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=2616;
					out<=216;
				end
				if(in == 3) begin
					state<=4516;
					out<=217;
				end
				if(in == 4) begin
					state<=618;
					out<=218;
				end
			end
			6495: begin
				if(in == 0) begin
					state<=6506;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=2617;
					out<=221;
				end
				if(in == 3) begin
					state<=4517;
					out<=222;
				end
				if(in == 4) begin
					state<=619;
					out<=223;
				end
			end
			6496: begin
				if(in == 0) begin
					state<=6507;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=2618;
					out<=226;
				end
				if(in == 3) begin
					state<=4518;
					out<=227;
				end
				if(in == 4) begin
					state<=620;
					out<=228;
				end
			end
			6497: begin
				if(in == 0) begin
					state<=6508;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=2619;
					out<=231;
				end
				if(in == 3) begin
					state<=4519;
					out<=232;
				end
				if(in == 4) begin
					state<=621;
					out<=233;
				end
			end
			6498: begin
				if(in == 0) begin
					state<=6499;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=2610;
					out<=236;
				end
				if(in == 3) begin
					state<=4510;
					out<=237;
				end
				if(in == 4) begin
					state<=612;
					out<=238;
				end
			end
			6499: begin
				if(in == 0) begin
					state<=6510;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=2621;
					out<=241;
				end
				if(in == 3) begin
					state<=4521;
					out<=242;
				end
				if(in == 4) begin
					state<=623;
					out<=243;
				end
			end
			6500: begin
				if(in == 0) begin
					state<=6511;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=2622;
					out<=246;
				end
				if(in == 3) begin
					state<=4522;
					out<=247;
				end
				if(in == 4) begin
					state<=624;
					out<=248;
				end
			end
			6501: begin
				if(in == 0) begin
					state<=6512;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=2623;
					out<=251;
				end
				if(in == 3) begin
					state<=4523;
					out<=252;
				end
				if(in == 4) begin
					state<=625;
					out<=253;
				end
			end
			6502: begin
				if(in == 0) begin
					state<=6513;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=2624;
					out<=0;
				end
				if(in == 3) begin
					state<=4524;
					out<=1;
				end
				if(in == 4) begin
					state<=626;
					out<=2;
				end
			end
			6503: begin
				if(in == 0) begin
					state<=6514;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=2625;
					out<=5;
				end
				if(in == 3) begin
					state<=4525;
					out<=6;
				end
				if(in == 4) begin
					state<=627;
					out<=7;
				end
			end
			6504: begin
				if(in == 0) begin
					state<=6515;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=2626;
					out<=10;
				end
				if(in == 3) begin
					state<=4526;
					out<=11;
				end
				if(in == 4) begin
					state<=628;
					out<=12;
				end
			end
			6505: begin
				if(in == 0) begin
					state<=6516;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=2627;
					out<=15;
				end
				if(in == 3) begin
					state<=4527;
					out<=16;
				end
				if(in == 4) begin
					state<=629;
					out<=17;
				end
			end
			6506: begin
				if(in == 0) begin
					state<=6517;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=2628;
					out<=20;
				end
				if(in == 3) begin
					state<=4528;
					out<=21;
				end
				if(in == 4) begin
					state<=630;
					out<=22;
				end
			end
			6507: begin
				if(in == 0) begin
					state<=6518;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=2629;
					out<=25;
				end
				if(in == 3) begin
					state<=4529;
					out<=26;
				end
				if(in == 4) begin
					state<=631;
					out<=27;
				end
			end
			6508: begin
				if(in == 0) begin
					state<=6509;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=2620;
					out<=30;
				end
				if(in == 3) begin
					state<=4520;
					out<=31;
				end
				if(in == 4) begin
					state<=622;
					out<=32;
				end
			end
			6509: begin
				if(in == 0) begin
					state<=6520;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=2631;
					out<=35;
				end
				if(in == 3) begin
					state<=4531;
					out<=36;
				end
				if(in == 4) begin
					state<=633;
					out<=37;
				end
			end
			6510: begin
				if(in == 0) begin
					state<=6521;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=2632;
					out<=40;
				end
				if(in == 3) begin
					state<=4532;
					out<=41;
				end
				if(in == 4) begin
					state<=634;
					out<=42;
				end
			end
			6511: begin
				if(in == 0) begin
					state<=6522;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=2633;
					out<=45;
				end
				if(in == 3) begin
					state<=4533;
					out<=46;
				end
				if(in == 4) begin
					state<=635;
					out<=47;
				end
			end
			6512: begin
				if(in == 0) begin
					state<=6523;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=2634;
					out<=50;
				end
				if(in == 3) begin
					state<=4534;
					out<=51;
				end
				if(in == 4) begin
					state<=636;
					out<=52;
				end
			end
			6513: begin
				if(in == 0) begin
					state<=6524;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=2635;
					out<=55;
				end
				if(in == 3) begin
					state<=4535;
					out<=56;
				end
				if(in == 4) begin
					state<=637;
					out<=57;
				end
			end
			6514: begin
				if(in == 0) begin
					state<=6525;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=2636;
					out<=60;
				end
				if(in == 3) begin
					state<=4536;
					out<=61;
				end
				if(in == 4) begin
					state<=638;
					out<=62;
				end
			end
			6515: begin
				if(in == 0) begin
					state<=6526;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=2637;
					out<=65;
				end
				if(in == 3) begin
					state<=4537;
					out<=66;
				end
				if(in == 4) begin
					state<=639;
					out<=67;
				end
			end
			6516: begin
				if(in == 0) begin
					state<=6527;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=2638;
					out<=70;
				end
				if(in == 3) begin
					state<=4538;
					out<=71;
				end
				if(in == 4) begin
					state<=640;
					out<=72;
				end
			end
			6517: begin
				if(in == 0) begin
					state<=6528;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=2639;
					out<=75;
				end
				if(in == 3) begin
					state<=4539;
					out<=76;
				end
				if(in == 4) begin
					state<=641;
					out<=77;
				end
			end
			6518: begin
				if(in == 0) begin
					state<=6519;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=2630;
					out<=80;
				end
				if(in == 3) begin
					state<=4530;
					out<=81;
				end
				if(in == 4) begin
					state<=632;
					out<=82;
				end
			end
			6519: begin
				if(in == 0) begin
					state<=6530;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=2641;
					out<=85;
				end
				if(in == 3) begin
					state<=4541;
					out<=86;
				end
				if(in == 4) begin
					state<=643;
					out<=87;
				end
			end
			6520: begin
				if(in == 0) begin
					state<=6531;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=2642;
					out<=90;
				end
				if(in == 3) begin
					state<=4542;
					out<=91;
				end
				if(in == 4) begin
					state<=644;
					out<=92;
				end
			end
			6521: begin
				if(in == 0) begin
					state<=6532;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=2643;
					out<=95;
				end
				if(in == 3) begin
					state<=4543;
					out<=96;
				end
				if(in == 4) begin
					state<=645;
					out<=97;
				end
			end
			6522: begin
				if(in == 0) begin
					state<=6533;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=2644;
					out<=100;
				end
				if(in == 3) begin
					state<=4544;
					out<=101;
				end
				if(in == 4) begin
					state<=646;
					out<=102;
				end
			end
			6523: begin
				if(in == 0) begin
					state<=6534;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=2645;
					out<=105;
				end
				if(in == 3) begin
					state<=4545;
					out<=106;
				end
				if(in == 4) begin
					state<=647;
					out<=107;
				end
			end
			6524: begin
				if(in == 0) begin
					state<=6535;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=2646;
					out<=110;
				end
				if(in == 3) begin
					state<=4546;
					out<=111;
				end
				if(in == 4) begin
					state<=648;
					out<=112;
				end
			end
			6525: begin
				if(in == 0) begin
					state<=6536;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=2647;
					out<=115;
				end
				if(in == 3) begin
					state<=4547;
					out<=116;
				end
				if(in == 4) begin
					state<=649;
					out<=117;
				end
			end
			6526: begin
				if(in == 0) begin
					state<=6537;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=2648;
					out<=120;
				end
				if(in == 3) begin
					state<=4548;
					out<=121;
				end
				if(in == 4) begin
					state<=650;
					out<=122;
				end
			end
			6527: begin
				if(in == 0) begin
					state<=6538;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=2649;
					out<=125;
				end
				if(in == 3) begin
					state<=4549;
					out<=126;
				end
				if(in == 4) begin
					state<=651;
					out<=127;
				end
			end
			6528: begin
				if(in == 0) begin
					state<=6529;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=2640;
					out<=130;
				end
				if(in == 3) begin
					state<=4540;
					out<=131;
				end
				if(in == 4) begin
					state<=642;
					out<=132;
				end
			end
			6529: begin
				if(in == 0) begin
					state<=6540;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=2651;
					out<=135;
				end
				if(in == 3) begin
					state<=4551;
					out<=136;
				end
				if(in == 4) begin
					state<=653;
					out<=137;
				end
			end
			6530: begin
				if(in == 0) begin
					state<=6541;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=2652;
					out<=140;
				end
				if(in == 3) begin
					state<=4552;
					out<=141;
				end
				if(in == 4) begin
					state<=654;
					out<=142;
				end
			end
			6531: begin
				if(in == 0) begin
					state<=6542;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=2653;
					out<=145;
				end
				if(in == 3) begin
					state<=4553;
					out<=146;
				end
				if(in == 4) begin
					state<=655;
					out<=147;
				end
			end
			6532: begin
				if(in == 0) begin
					state<=6543;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=2654;
					out<=150;
				end
				if(in == 3) begin
					state<=4554;
					out<=151;
				end
				if(in == 4) begin
					state<=656;
					out<=152;
				end
			end
			6533: begin
				if(in == 0) begin
					state<=6544;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=2655;
					out<=155;
				end
				if(in == 3) begin
					state<=4555;
					out<=156;
				end
				if(in == 4) begin
					state<=657;
					out<=157;
				end
			end
			6534: begin
				if(in == 0) begin
					state<=6545;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=2656;
					out<=160;
				end
				if(in == 3) begin
					state<=4556;
					out<=161;
				end
				if(in == 4) begin
					state<=658;
					out<=162;
				end
			end
			6535: begin
				if(in == 0) begin
					state<=6546;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=2657;
					out<=165;
				end
				if(in == 3) begin
					state<=4557;
					out<=166;
				end
				if(in == 4) begin
					state<=659;
					out<=167;
				end
			end
			6536: begin
				if(in == 0) begin
					state<=6547;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=2658;
					out<=170;
				end
				if(in == 3) begin
					state<=4558;
					out<=171;
				end
				if(in == 4) begin
					state<=660;
					out<=172;
				end
			end
			6537: begin
				if(in == 0) begin
					state<=6548;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=2659;
					out<=175;
				end
				if(in == 3) begin
					state<=4559;
					out<=176;
				end
				if(in == 4) begin
					state<=661;
					out<=177;
				end
			end
			6538: begin
				if(in == 0) begin
					state<=6539;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=2650;
					out<=180;
				end
				if(in == 3) begin
					state<=4550;
					out<=181;
				end
				if(in == 4) begin
					state<=652;
					out<=182;
				end
			end
			6539: begin
				if(in == 0) begin
					state<=6550;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=2661;
					out<=185;
				end
				if(in == 3) begin
					state<=4561;
					out<=186;
				end
				if(in == 4) begin
					state<=663;
					out<=187;
				end
			end
			6540: begin
				if(in == 0) begin
					state<=6551;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=2662;
					out<=190;
				end
				if(in == 3) begin
					state<=4562;
					out<=191;
				end
				if(in == 4) begin
					state<=664;
					out<=192;
				end
			end
			6541: begin
				if(in == 0) begin
					state<=6552;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=2663;
					out<=195;
				end
				if(in == 3) begin
					state<=4563;
					out<=196;
				end
				if(in == 4) begin
					state<=665;
					out<=197;
				end
			end
			6542: begin
				if(in == 0) begin
					state<=6553;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=2664;
					out<=200;
				end
				if(in == 3) begin
					state<=4564;
					out<=201;
				end
				if(in == 4) begin
					state<=666;
					out<=202;
				end
			end
			6543: begin
				if(in == 0) begin
					state<=6554;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=2665;
					out<=205;
				end
				if(in == 3) begin
					state<=4565;
					out<=206;
				end
				if(in == 4) begin
					state<=667;
					out<=207;
				end
			end
			6544: begin
				if(in == 0) begin
					state<=6555;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=2666;
					out<=210;
				end
				if(in == 3) begin
					state<=4566;
					out<=211;
				end
				if(in == 4) begin
					state<=668;
					out<=212;
				end
			end
			6545: begin
				if(in == 0) begin
					state<=6556;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=2667;
					out<=215;
				end
				if(in == 3) begin
					state<=4567;
					out<=216;
				end
				if(in == 4) begin
					state<=669;
					out<=217;
				end
			end
			6546: begin
				if(in == 0) begin
					state<=6557;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=2668;
					out<=220;
				end
				if(in == 3) begin
					state<=4568;
					out<=221;
				end
				if(in == 4) begin
					state<=670;
					out<=222;
				end
			end
			6547: begin
				if(in == 0) begin
					state<=6558;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=2669;
					out<=225;
				end
				if(in == 3) begin
					state<=4569;
					out<=226;
				end
				if(in == 4) begin
					state<=671;
					out<=227;
				end
			end
			6548: begin
				if(in == 0) begin
					state<=6549;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=2660;
					out<=230;
				end
				if(in == 3) begin
					state<=4560;
					out<=231;
				end
				if(in == 4) begin
					state<=662;
					out<=232;
				end
			end
			6549: begin
				if(in == 0) begin
					state<=7120;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=3231;
					out<=235;
				end
				if(in == 3) begin
					state<=5467;
					out<=236;
				end
				if(in == 4) begin
					state<=1578;
					out<=237;
				end
			end
			6550: begin
				if(in == 0) begin
					state<=7121;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=3232;
					out<=240;
				end
				if(in == 3) begin
					state<=5468;
					out<=241;
				end
				if(in == 4) begin
					state<=1579;
					out<=242;
				end
			end
			6551: begin
				if(in == 0) begin
					state<=7122;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=3233;
					out<=245;
				end
				if(in == 3) begin
					state<=5469;
					out<=246;
				end
				if(in == 4) begin
					state<=1580;
					out<=247;
				end
			end
			6552: begin
				if(in == 0) begin
					state<=7123;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=3234;
					out<=250;
				end
				if(in == 3) begin
					state<=5470;
					out<=251;
				end
				if(in == 4) begin
					state<=1581;
					out<=252;
				end
			end
			6553: begin
				if(in == 0) begin
					state<=7124;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=3235;
					out<=255;
				end
				if(in == 3) begin
					state<=5471;
					out<=0;
				end
				if(in == 4) begin
					state<=1582;
					out<=1;
				end
			end
			6554: begin
				if(in == 0) begin
					state<=7125;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=3236;
					out<=4;
				end
				if(in == 3) begin
					state<=5472;
					out<=5;
				end
				if(in == 4) begin
					state<=1583;
					out<=6;
				end
			end
			6555: begin
				if(in == 0) begin
					state<=7126;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=3237;
					out<=9;
				end
				if(in == 3) begin
					state<=5473;
					out<=10;
				end
				if(in == 4) begin
					state<=1584;
					out<=11;
				end
			end
			6556: begin
				if(in == 0) begin
					state<=7127;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=3238;
					out<=14;
				end
				if(in == 3) begin
					state<=5474;
					out<=15;
				end
				if(in == 4) begin
					state<=1585;
					out<=16;
				end
			end
			6557: begin
				if(in == 0) begin
					state<=7128;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=3239;
					out<=19;
				end
				if(in == 3) begin
					state<=5475;
					out<=20;
				end
				if(in == 4) begin
					state<=1586;
					out<=21;
				end
			end
			6558: begin
				if(in == 0) begin
					state<=7119;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=3230;
					out<=24;
				end
				if(in == 3) begin
					state<=5466;
					out<=25;
				end
				if(in == 4) begin
					state<=1577;
					out<=26;
				end
			end
			6559: begin
				if(in == 0) begin
					state<=6570;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=2681;
					out<=29;
				end
				if(in == 3) begin
					state<=4581;
					out<=30;
				end
				if(in == 4) begin
					state<=683;
					out<=31;
				end
			end
			6560: begin
				if(in == 0) begin
					state<=6571;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=2682;
					out<=34;
				end
				if(in == 3) begin
					state<=4582;
					out<=35;
				end
				if(in == 4) begin
					state<=684;
					out<=36;
				end
			end
			6561: begin
				if(in == 0) begin
					state<=6572;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=2683;
					out<=39;
				end
				if(in == 3) begin
					state<=4583;
					out<=40;
				end
				if(in == 4) begin
					state<=685;
					out<=41;
				end
			end
			6562: begin
				if(in == 0) begin
					state<=6573;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=2684;
					out<=44;
				end
				if(in == 3) begin
					state<=4584;
					out<=45;
				end
				if(in == 4) begin
					state<=686;
					out<=46;
				end
			end
			6563: begin
				if(in == 0) begin
					state<=6574;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=2685;
					out<=49;
				end
				if(in == 3) begin
					state<=4585;
					out<=50;
				end
				if(in == 4) begin
					state<=687;
					out<=51;
				end
			end
			6564: begin
				if(in == 0) begin
					state<=6575;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=2686;
					out<=54;
				end
				if(in == 3) begin
					state<=4586;
					out<=55;
				end
				if(in == 4) begin
					state<=688;
					out<=56;
				end
			end
			6565: begin
				if(in == 0) begin
					state<=6576;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=2687;
					out<=59;
				end
				if(in == 3) begin
					state<=4587;
					out<=60;
				end
				if(in == 4) begin
					state<=689;
					out<=61;
				end
			end
			6566: begin
				if(in == 0) begin
					state<=6577;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=2688;
					out<=64;
				end
				if(in == 3) begin
					state<=4588;
					out<=65;
				end
				if(in == 4) begin
					state<=690;
					out<=66;
				end
			end
			6567: begin
				if(in == 0) begin
					state<=6568;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=2679;
					out<=69;
				end
				if(in == 3) begin
					state<=4579;
					out<=70;
				end
				if(in == 4) begin
					state<=681;
					out<=71;
				end
			end
			6568: begin
				if(in == 0) begin
					state<=5889;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=2000;
					out<=74;
				end
				if(in == 3) begin
					state<=3900;
					out<=75;
				end
				if(in == 4) begin
					state<=2;
					out<=76;
				end
			end
			6569: begin
				if(in == 0) begin
					state<=5890;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=2001;
					out<=79;
				end
				if(in == 3) begin
					state<=3901;
					out<=80;
				end
				if(in == 4) begin
					state<=3;
					out<=81;
				end
			end
			6570: begin
				if(in == 0) begin
					state<=5891;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=2002;
					out<=84;
				end
				if(in == 3) begin
					state<=3902;
					out<=85;
				end
				if(in == 4) begin
					state<=4;
					out<=86;
				end
			end
			6571: begin
				if(in == 0) begin
					state<=5892;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=2003;
					out<=89;
				end
				if(in == 3) begin
					state<=3903;
					out<=90;
				end
				if(in == 4) begin
					state<=5;
					out<=91;
				end
			end
			6572: begin
				if(in == 0) begin
					state<=5893;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=2004;
					out<=94;
				end
				if(in == 3) begin
					state<=3904;
					out<=95;
				end
				if(in == 4) begin
					state<=6;
					out<=96;
				end
			end
			6573: begin
				if(in == 0) begin
					state<=5894;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=2005;
					out<=99;
				end
				if(in == 3) begin
					state<=3905;
					out<=100;
				end
				if(in == 4) begin
					state<=7;
					out<=101;
				end
			end
			6574: begin
				if(in == 0) begin
					state<=5895;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=2006;
					out<=104;
				end
				if(in == 3) begin
					state<=3906;
					out<=105;
				end
				if(in == 4) begin
					state<=8;
					out<=106;
				end
			end
			6575: begin
				if(in == 0) begin
					state<=5896;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=2007;
					out<=109;
				end
				if(in == 3) begin
					state<=3907;
					out<=110;
				end
				if(in == 4) begin
					state<=9;
					out<=111;
				end
			end
			6576: begin
				if(in == 0) begin
					state<=5897;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=2008;
					out<=114;
				end
				if(in == 3) begin
					state<=3908;
					out<=115;
				end
				if(in == 4) begin
					state<=10;
					out<=116;
				end
			end
			6577: begin
				if(in == 0) begin
					state<=5888;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=1999;
					out<=119;
				end
				if(in == 3) begin
					state<=3899;
					out<=120;
				end
				if(in == 4) begin
					state<=1;
					out<=121;
				end
			end
			6578: begin
				if(in == 0) begin
					state<=6589;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=2700;
					out<=124;
				end
				if(in == 3) begin
					state<=4600;
					out<=125;
				end
				if(in == 4) begin
					state<=702;
					out<=126;
				end
			end
			6579: begin
				if(in == 0) begin
					state<=6590;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=2701;
					out<=129;
				end
				if(in == 3) begin
					state<=4601;
					out<=130;
				end
				if(in == 4) begin
					state<=703;
					out<=131;
				end
			end
			6580: begin
				if(in == 0) begin
					state<=6591;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=2702;
					out<=134;
				end
				if(in == 3) begin
					state<=4602;
					out<=135;
				end
				if(in == 4) begin
					state<=704;
					out<=136;
				end
			end
			6581: begin
				if(in == 0) begin
					state<=6592;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=2703;
					out<=139;
				end
				if(in == 3) begin
					state<=4603;
					out<=140;
				end
				if(in == 4) begin
					state<=705;
					out<=141;
				end
			end
			6582: begin
				if(in == 0) begin
					state<=6593;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=2704;
					out<=144;
				end
				if(in == 3) begin
					state<=4604;
					out<=145;
				end
				if(in == 4) begin
					state<=706;
					out<=146;
				end
			end
			6583: begin
				if(in == 0) begin
					state<=6594;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=2705;
					out<=149;
				end
				if(in == 3) begin
					state<=4605;
					out<=150;
				end
				if(in == 4) begin
					state<=707;
					out<=151;
				end
			end
			6584: begin
				if(in == 0) begin
					state<=6595;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=2706;
					out<=154;
				end
				if(in == 3) begin
					state<=4606;
					out<=155;
				end
				if(in == 4) begin
					state<=708;
					out<=156;
				end
			end
			6585: begin
				if(in == 0) begin
					state<=6596;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=2707;
					out<=159;
				end
				if(in == 3) begin
					state<=4607;
					out<=160;
				end
				if(in == 4) begin
					state<=709;
					out<=161;
				end
			end
			6586: begin
				if(in == 0) begin
					state<=6587;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=2698;
					out<=164;
				end
				if(in == 3) begin
					state<=4598;
					out<=165;
				end
				if(in == 4) begin
					state<=700;
					out<=166;
				end
			end
			6587: begin
				if(in == 0) begin
					state<=6598;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=2709;
					out<=169;
				end
				if(in == 3) begin
					state<=4609;
					out<=170;
				end
				if(in == 4) begin
					state<=711;
					out<=171;
				end
			end
			6588: begin
				if(in == 0) begin
					state<=6599;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=2710;
					out<=174;
				end
				if(in == 3) begin
					state<=4610;
					out<=175;
				end
				if(in == 4) begin
					state<=712;
					out<=176;
				end
			end
			6589: begin
				if(in == 0) begin
					state<=6600;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=2711;
					out<=179;
				end
				if(in == 3) begin
					state<=4611;
					out<=180;
				end
				if(in == 4) begin
					state<=713;
					out<=181;
				end
			end
			6590: begin
				if(in == 0) begin
					state<=6601;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=2712;
					out<=184;
				end
				if(in == 3) begin
					state<=4612;
					out<=185;
				end
				if(in == 4) begin
					state<=714;
					out<=186;
				end
			end
			6591: begin
				if(in == 0) begin
					state<=6602;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=2713;
					out<=189;
				end
				if(in == 3) begin
					state<=4613;
					out<=190;
				end
				if(in == 4) begin
					state<=715;
					out<=191;
				end
			end
			6592: begin
				if(in == 0) begin
					state<=6603;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=2714;
					out<=194;
				end
				if(in == 3) begin
					state<=4614;
					out<=195;
				end
				if(in == 4) begin
					state<=716;
					out<=196;
				end
			end
			6593: begin
				if(in == 0) begin
					state<=6604;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=2715;
					out<=199;
				end
				if(in == 3) begin
					state<=4615;
					out<=200;
				end
				if(in == 4) begin
					state<=717;
					out<=201;
				end
			end
			6594: begin
				if(in == 0) begin
					state<=6605;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=2716;
					out<=204;
				end
				if(in == 3) begin
					state<=4616;
					out<=205;
				end
				if(in == 4) begin
					state<=718;
					out<=206;
				end
			end
			6595: begin
				if(in == 0) begin
					state<=6606;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=2717;
					out<=209;
				end
				if(in == 3) begin
					state<=4617;
					out<=210;
				end
				if(in == 4) begin
					state<=719;
					out<=211;
				end
			end
			6596: begin
				if(in == 0) begin
					state<=6597;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=2708;
					out<=214;
				end
				if(in == 3) begin
					state<=4608;
					out<=215;
				end
				if(in == 4) begin
					state<=710;
					out<=216;
				end
			end
			6597: begin
				if(in == 0) begin
					state<=6608;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=2719;
					out<=219;
				end
				if(in == 3) begin
					state<=4619;
					out<=220;
				end
				if(in == 4) begin
					state<=721;
					out<=221;
				end
			end
			6598: begin
				if(in == 0) begin
					state<=6609;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=2720;
					out<=224;
				end
				if(in == 3) begin
					state<=4620;
					out<=225;
				end
				if(in == 4) begin
					state<=722;
					out<=226;
				end
			end
			6599: begin
				if(in == 0) begin
					state<=6610;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=2721;
					out<=229;
				end
				if(in == 3) begin
					state<=4621;
					out<=230;
				end
				if(in == 4) begin
					state<=723;
					out<=231;
				end
			end
			6600: begin
				if(in == 0) begin
					state<=6611;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=2722;
					out<=234;
				end
				if(in == 3) begin
					state<=4622;
					out<=235;
				end
				if(in == 4) begin
					state<=724;
					out<=236;
				end
			end
			6601: begin
				if(in == 0) begin
					state<=6612;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=2723;
					out<=239;
				end
				if(in == 3) begin
					state<=4623;
					out<=240;
				end
				if(in == 4) begin
					state<=725;
					out<=241;
				end
			end
			6602: begin
				if(in == 0) begin
					state<=6613;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=2724;
					out<=244;
				end
				if(in == 3) begin
					state<=4624;
					out<=245;
				end
				if(in == 4) begin
					state<=726;
					out<=246;
				end
			end
			6603: begin
				if(in == 0) begin
					state<=6614;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=2725;
					out<=249;
				end
				if(in == 3) begin
					state<=4625;
					out<=250;
				end
				if(in == 4) begin
					state<=727;
					out<=251;
				end
			end
			6604: begin
				if(in == 0) begin
					state<=6615;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=2726;
					out<=254;
				end
				if(in == 3) begin
					state<=4626;
					out<=255;
				end
				if(in == 4) begin
					state<=728;
					out<=0;
				end
			end
			6605: begin
				if(in == 0) begin
					state<=6616;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=2727;
					out<=3;
				end
				if(in == 3) begin
					state<=4627;
					out<=4;
				end
				if(in == 4) begin
					state<=729;
					out<=5;
				end
			end
			6606: begin
				if(in == 0) begin
					state<=6607;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=2718;
					out<=8;
				end
				if(in == 3) begin
					state<=4618;
					out<=9;
				end
				if(in == 4) begin
					state<=720;
					out<=10;
				end
			end
			6607: begin
				if(in == 0) begin
					state<=6618;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=2729;
					out<=13;
				end
				if(in == 3) begin
					state<=4629;
					out<=14;
				end
				if(in == 4) begin
					state<=731;
					out<=15;
				end
			end
			6608: begin
				if(in == 0) begin
					state<=6619;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=2730;
					out<=18;
				end
				if(in == 3) begin
					state<=4630;
					out<=19;
				end
				if(in == 4) begin
					state<=732;
					out<=20;
				end
			end
			6609: begin
				if(in == 0) begin
					state<=6620;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=2731;
					out<=23;
				end
				if(in == 3) begin
					state<=4631;
					out<=24;
				end
				if(in == 4) begin
					state<=733;
					out<=25;
				end
			end
			6610: begin
				if(in == 0) begin
					state<=6621;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=2732;
					out<=28;
				end
				if(in == 3) begin
					state<=4632;
					out<=29;
				end
				if(in == 4) begin
					state<=734;
					out<=30;
				end
			end
			6611: begin
				if(in == 0) begin
					state<=6622;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=2733;
					out<=33;
				end
				if(in == 3) begin
					state<=4633;
					out<=34;
				end
				if(in == 4) begin
					state<=735;
					out<=35;
				end
			end
			6612: begin
				if(in == 0) begin
					state<=6623;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=2734;
					out<=38;
				end
				if(in == 3) begin
					state<=4634;
					out<=39;
				end
				if(in == 4) begin
					state<=736;
					out<=40;
				end
			end
			6613: begin
				if(in == 0) begin
					state<=6624;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=2735;
					out<=43;
				end
				if(in == 3) begin
					state<=4635;
					out<=44;
				end
				if(in == 4) begin
					state<=737;
					out<=45;
				end
			end
			6614: begin
				if(in == 0) begin
					state<=6625;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=2736;
					out<=48;
				end
				if(in == 3) begin
					state<=4636;
					out<=49;
				end
				if(in == 4) begin
					state<=738;
					out<=50;
				end
			end
			6615: begin
				if(in == 0) begin
					state<=6626;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=2737;
					out<=53;
				end
				if(in == 3) begin
					state<=4637;
					out<=54;
				end
				if(in == 4) begin
					state<=739;
					out<=55;
				end
			end
			6616: begin
				if(in == 0) begin
					state<=6617;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=2728;
					out<=58;
				end
				if(in == 3) begin
					state<=4628;
					out<=59;
				end
				if(in == 4) begin
					state<=730;
					out<=60;
				end
			end
			6617: begin
				if(in == 0) begin
					state<=6628;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=2739;
					out<=63;
				end
				if(in == 3) begin
					state<=4639;
					out<=64;
				end
				if(in == 4) begin
					state<=741;
					out<=65;
				end
			end
			6618: begin
				if(in == 0) begin
					state<=6629;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=2740;
					out<=68;
				end
				if(in == 3) begin
					state<=4640;
					out<=69;
				end
				if(in == 4) begin
					state<=742;
					out<=70;
				end
			end
			6619: begin
				if(in == 0) begin
					state<=6630;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=2741;
					out<=73;
				end
				if(in == 3) begin
					state<=4641;
					out<=74;
				end
				if(in == 4) begin
					state<=743;
					out<=75;
				end
			end
			6620: begin
				if(in == 0) begin
					state<=6631;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=2742;
					out<=78;
				end
				if(in == 3) begin
					state<=4642;
					out<=79;
				end
				if(in == 4) begin
					state<=744;
					out<=80;
				end
			end
			6621: begin
				if(in == 0) begin
					state<=6632;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=2743;
					out<=83;
				end
				if(in == 3) begin
					state<=4643;
					out<=84;
				end
				if(in == 4) begin
					state<=745;
					out<=85;
				end
			end
			6622: begin
				if(in == 0) begin
					state<=6633;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=2744;
					out<=88;
				end
				if(in == 3) begin
					state<=4644;
					out<=89;
				end
				if(in == 4) begin
					state<=746;
					out<=90;
				end
			end
			6623: begin
				if(in == 0) begin
					state<=6634;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=2745;
					out<=93;
				end
				if(in == 3) begin
					state<=4645;
					out<=94;
				end
				if(in == 4) begin
					state<=747;
					out<=95;
				end
			end
			6624: begin
				if(in == 0) begin
					state<=6635;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=2746;
					out<=98;
				end
				if(in == 3) begin
					state<=4646;
					out<=99;
				end
				if(in == 4) begin
					state<=748;
					out<=100;
				end
			end
			6625: begin
				if(in == 0) begin
					state<=6636;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=2747;
					out<=103;
				end
				if(in == 3) begin
					state<=4647;
					out<=104;
				end
				if(in == 4) begin
					state<=749;
					out<=105;
				end
			end
			6626: begin
				if(in == 0) begin
					state<=6627;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=2738;
					out<=108;
				end
				if(in == 3) begin
					state<=4638;
					out<=109;
				end
				if(in == 4) begin
					state<=740;
					out<=110;
				end
			end
			6627: begin
				if(in == 0) begin
					state<=6638;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=2749;
					out<=113;
				end
				if(in == 3) begin
					state<=4649;
					out<=114;
				end
				if(in == 4) begin
					state<=751;
					out<=115;
				end
			end
			6628: begin
				if(in == 0) begin
					state<=6639;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=2750;
					out<=118;
				end
				if(in == 3) begin
					state<=4650;
					out<=119;
				end
				if(in == 4) begin
					state<=752;
					out<=120;
				end
			end
			6629: begin
				if(in == 0) begin
					state<=6640;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=2751;
					out<=123;
				end
				if(in == 3) begin
					state<=4651;
					out<=124;
				end
				if(in == 4) begin
					state<=753;
					out<=125;
				end
			end
			6630: begin
				if(in == 0) begin
					state<=6641;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=2752;
					out<=128;
				end
				if(in == 3) begin
					state<=4652;
					out<=129;
				end
				if(in == 4) begin
					state<=754;
					out<=130;
				end
			end
			6631: begin
				if(in == 0) begin
					state<=6642;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=2753;
					out<=133;
				end
				if(in == 3) begin
					state<=4653;
					out<=134;
				end
				if(in == 4) begin
					state<=755;
					out<=135;
				end
			end
			6632: begin
				if(in == 0) begin
					state<=6643;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=2754;
					out<=138;
				end
				if(in == 3) begin
					state<=4654;
					out<=139;
				end
				if(in == 4) begin
					state<=756;
					out<=140;
				end
			end
			6633: begin
				if(in == 0) begin
					state<=6644;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=2755;
					out<=143;
				end
				if(in == 3) begin
					state<=4655;
					out<=144;
				end
				if(in == 4) begin
					state<=757;
					out<=145;
				end
			end
			6634: begin
				if(in == 0) begin
					state<=6645;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=2756;
					out<=148;
				end
				if(in == 3) begin
					state<=4656;
					out<=149;
				end
				if(in == 4) begin
					state<=758;
					out<=150;
				end
			end
			6635: begin
				if(in == 0) begin
					state<=6646;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=2757;
					out<=153;
				end
				if(in == 3) begin
					state<=4657;
					out<=154;
				end
				if(in == 4) begin
					state<=759;
					out<=155;
				end
			end
			6636: begin
				if(in == 0) begin
					state<=6637;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=2748;
					out<=158;
				end
				if(in == 3) begin
					state<=4648;
					out<=159;
				end
				if(in == 4) begin
					state<=750;
					out<=160;
				end
			end
			6637: begin
				if(in == 0) begin
					state<=6648;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=2759;
					out<=163;
				end
				if(in == 3) begin
					state<=4659;
					out<=164;
				end
				if(in == 4) begin
					state<=761;
					out<=165;
				end
			end
			6638: begin
				if(in == 0) begin
					state<=6649;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=2760;
					out<=168;
				end
				if(in == 3) begin
					state<=4660;
					out<=169;
				end
				if(in == 4) begin
					state<=762;
					out<=170;
				end
			end
			6639: begin
				if(in == 0) begin
					state<=6650;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=2761;
					out<=173;
				end
				if(in == 3) begin
					state<=4661;
					out<=174;
				end
				if(in == 4) begin
					state<=763;
					out<=175;
				end
			end
			6640: begin
				if(in == 0) begin
					state<=6651;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=2762;
					out<=178;
				end
				if(in == 3) begin
					state<=4662;
					out<=179;
				end
				if(in == 4) begin
					state<=764;
					out<=180;
				end
			end
			6641: begin
				if(in == 0) begin
					state<=6652;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=2763;
					out<=183;
				end
				if(in == 3) begin
					state<=4663;
					out<=184;
				end
				if(in == 4) begin
					state<=765;
					out<=185;
				end
			end
			6642: begin
				if(in == 0) begin
					state<=6653;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=2764;
					out<=188;
				end
				if(in == 3) begin
					state<=4664;
					out<=189;
				end
				if(in == 4) begin
					state<=766;
					out<=190;
				end
			end
			6643: begin
				if(in == 0) begin
					state<=6654;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=2765;
					out<=193;
				end
				if(in == 3) begin
					state<=4665;
					out<=194;
				end
				if(in == 4) begin
					state<=767;
					out<=195;
				end
			end
			6644: begin
				if(in == 0) begin
					state<=6655;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=2766;
					out<=198;
				end
				if(in == 3) begin
					state<=4666;
					out<=199;
				end
				if(in == 4) begin
					state<=768;
					out<=200;
				end
			end
			6645: begin
				if(in == 0) begin
					state<=6656;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=2767;
					out<=203;
				end
				if(in == 3) begin
					state<=4667;
					out<=204;
				end
				if(in == 4) begin
					state<=769;
					out<=205;
				end
			end
			6646: begin
				if(in == 0) begin
					state<=6647;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=2758;
					out<=208;
				end
				if(in == 3) begin
					state<=4658;
					out<=209;
				end
				if(in == 4) begin
					state<=760;
					out<=210;
				end
			end
			6647: begin
				if(in == 0) begin
					state<=6658;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=2769;
					out<=213;
				end
				if(in == 3) begin
					state<=4669;
					out<=214;
				end
				if(in == 4) begin
					state<=771;
					out<=215;
				end
			end
			6648: begin
				if(in == 0) begin
					state<=6659;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=2770;
					out<=218;
				end
				if(in == 3) begin
					state<=4670;
					out<=219;
				end
				if(in == 4) begin
					state<=772;
					out<=220;
				end
			end
			6649: begin
				if(in == 0) begin
					state<=6660;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=2771;
					out<=223;
				end
				if(in == 3) begin
					state<=4671;
					out<=224;
				end
				if(in == 4) begin
					state<=773;
					out<=225;
				end
			end
			6650: begin
				if(in == 0) begin
					state<=6661;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=2772;
					out<=228;
				end
				if(in == 3) begin
					state<=4672;
					out<=229;
				end
				if(in == 4) begin
					state<=774;
					out<=230;
				end
			end
			6651: begin
				if(in == 0) begin
					state<=6662;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=2773;
					out<=233;
				end
				if(in == 3) begin
					state<=4673;
					out<=234;
				end
				if(in == 4) begin
					state<=775;
					out<=235;
				end
			end
			6652: begin
				if(in == 0) begin
					state<=6663;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=2774;
					out<=238;
				end
				if(in == 3) begin
					state<=4674;
					out<=239;
				end
				if(in == 4) begin
					state<=776;
					out<=240;
				end
			end
			6653: begin
				if(in == 0) begin
					state<=6664;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=2775;
					out<=243;
				end
				if(in == 3) begin
					state<=4675;
					out<=244;
				end
				if(in == 4) begin
					state<=777;
					out<=245;
				end
			end
			6654: begin
				if(in == 0) begin
					state<=6665;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=2776;
					out<=248;
				end
				if(in == 3) begin
					state<=4676;
					out<=249;
				end
				if(in == 4) begin
					state<=778;
					out<=250;
				end
			end
			6655: begin
				if(in == 0) begin
					state<=6666;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=2777;
					out<=253;
				end
				if(in == 3) begin
					state<=4677;
					out<=254;
				end
				if(in == 4) begin
					state<=779;
					out<=255;
				end
			end
			6656: begin
				if(in == 0) begin
					state<=6657;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=2768;
					out<=2;
				end
				if(in == 3) begin
					state<=4668;
					out<=3;
				end
				if(in == 4) begin
					state<=770;
					out<=4;
				end
			end
			6657: begin
				if(in == 0) begin
					state<=6668;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=2779;
					out<=7;
				end
				if(in == 3) begin
					state<=4679;
					out<=8;
				end
				if(in == 4) begin
					state<=781;
					out<=9;
				end
			end
			6658: begin
				if(in == 0) begin
					state<=6669;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=2780;
					out<=12;
				end
				if(in == 3) begin
					state<=4680;
					out<=13;
				end
				if(in == 4) begin
					state<=782;
					out<=14;
				end
			end
			6659: begin
				if(in == 0) begin
					state<=6670;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=2781;
					out<=17;
				end
				if(in == 3) begin
					state<=4681;
					out<=18;
				end
				if(in == 4) begin
					state<=783;
					out<=19;
				end
			end
			6660: begin
				if(in == 0) begin
					state<=6671;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=2782;
					out<=22;
				end
				if(in == 3) begin
					state<=4682;
					out<=23;
				end
				if(in == 4) begin
					state<=784;
					out<=24;
				end
			end
			6661: begin
				if(in == 0) begin
					state<=6672;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=2783;
					out<=27;
				end
				if(in == 3) begin
					state<=4683;
					out<=28;
				end
				if(in == 4) begin
					state<=785;
					out<=29;
				end
			end
			6662: begin
				if(in == 0) begin
					state<=6673;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=2784;
					out<=32;
				end
				if(in == 3) begin
					state<=4684;
					out<=33;
				end
				if(in == 4) begin
					state<=786;
					out<=34;
				end
			end
			6663: begin
				if(in == 0) begin
					state<=6674;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=2785;
					out<=37;
				end
				if(in == 3) begin
					state<=4685;
					out<=38;
				end
				if(in == 4) begin
					state<=787;
					out<=39;
				end
			end
			6664: begin
				if(in == 0) begin
					state<=6675;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=2786;
					out<=42;
				end
				if(in == 3) begin
					state<=4686;
					out<=43;
				end
				if(in == 4) begin
					state<=788;
					out<=44;
				end
			end
			6665: begin
				if(in == 0) begin
					state<=6676;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=2787;
					out<=47;
				end
				if(in == 3) begin
					state<=4687;
					out<=48;
				end
				if(in == 4) begin
					state<=789;
					out<=49;
				end
			end
			6666: begin
				if(in == 0) begin
					state<=6667;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=2778;
					out<=52;
				end
				if(in == 3) begin
					state<=4678;
					out<=53;
				end
				if(in == 4) begin
					state<=780;
					out<=54;
				end
			end
			6667: begin
				if(in == 0) begin
					state<=6678;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=2789;
					out<=57;
				end
				if(in == 3) begin
					state<=4689;
					out<=58;
				end
				if(in == 4) begin
					state<=791;
					out<=59;
				end
			end
			6668: begin
				if(in == 0) begin
					state<=6679;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=2790;
					out<=62;
				end
				if(in == 3) begin
					state<=4690;
					out<=63;
				end
				if(in == 4) begin
					state<=792;
					out<=64;
				end
			end
			6669: begin
				if(in == 0) begin
					state<=6680;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=2791;
					out<=67;
				end
				if(in == 3) begin
					state<=4691;
					out<=68;
				end
				if(in == 4) begin
					state<=793;
					out<=69;
				end
			end
			6670: begin
				if(in == 0) begin
					state<=6681;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=2792;
					out<=72;
				end
				if(in == 3) begin
					state<=4692;
					out<=73;
				end
				if(in == 4) begin
					state<=794;
					out<=74;
				end
			end
			6671: begin
				if(in == 0) begin
					state<=6682;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=2793;
					out<=77;
				end
				if(in == 3) begin
					state<=4693;
					out<=78;
				end
				if(in == 4) begin
					state<=795;
					out<=79;
				end
			end
			6672: begin
				if(in == 0) begin
					state<=6683;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=2794;
					out<=82;
				end
				if(in == 3) begin
					state<=4694;
					out<=83;
				end
				if(in == 4) begin
					state<=796;
					out<=84;
				end
			end
			6673: begin
				if(in == 0) begin
					state<=6684;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=2795;
					out<=87;
				end
				if(in == 3) begin
					state<=4695;
					out<=88;
				end
				if(in == 4) begin
					state<=797;
					out<=89;
				end
			end
			6674: begin
				if(in == 0) begin
					state<=6685;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=2796;
					out<=92;
				end
				if(in == 3) begin
					state<=4696;
					out<=93;
				end
				if(in == 4) begin
					state<=798;
					out<=94;
				end
			end
			6675: begin
				if(in == 0) begin
					state<=6686;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=2797;
					out<=97;
				end
				if(in == 3) begin
					state<=4697;
					out<=98;
				end
				if(in == 4) begin
					state<=799;
					out<=99;
				end
			end
			6676: begin
				if(in == 0) begin
					state<=6677;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=2788;
					out<=102;
				end
				if(in == 3) begin
					state<=4688;
					out<=103;
				end
				if(in == 4) begin
					state<=790;
					out<=104;
				end
			end
			6677: begin
				if(in == 0) begin
					state<=6698;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=2809;
					out<=107;
				end
				if(in == 3) begin
					state<=4709;
					out<=108;
				end
				if(in == 4) begin
					state<=811;
					out<=109;
				end
			end
			6678: begin
				if(in == 0) begin
					state<=6699;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=2810;
					out<=112;
				end
				if(in == 3) begin
					state<=4710;
					out<=113;
				end
				if(in == 4) begin
					state<=812;
					out<=114;
				end
			end
			6679: begin
				if(in == 0) begin
					state<=6700;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=2811;
					out<=117;
				end
				if(in == 3) begin
					state<=4711;
					out<=118;
				end
				if(in == 4) begin
					state<=813;
					out<=119;
				end
			end
			6680: begin
				if(in == 0) begin
					state<=6701;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=2812;
					out<=122;
				end
				if(in == 3) begin
					state<=4712;
					out<=123;
				end
				if(in == 4) begin
					state<=814;
					out<=124;
				end
			end
			6681: begin
				if(in == 0) begin
					state<=6702;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=2813;
					out<=127;
				end
				if(in == 3) begin
					state<=4713;
					out<=128;
				end
				if(in == 4) begin
					state<=815;
					out<=129;
				end
			end
			6682: begin
				if(in == 0) begin
					state<=6703;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=2814;
					out<=132;
				end
				if(in == 3) begin
					state<=4714;
					out<=133;
				end
				if(in == 4) begin
					state<=816;
					out<=134;
				end
			end
			6683: begin
				if(in == 0) begin
					state<=6704;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=2815;
					out<=137;
				end
				if(in == 3) begin
					state<=4715;
					out<=138;
				end
				if(in == 4) begin
					state<=817;
					out<=139;
				end
			end
			6684: begin
				if(in == 0) begin
					state<=6705;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=2816;
					out<=142;
				end
				if(in == 3) begin
					state<=4716;
					out<=143;
				end
				if(in == 4) begin
					state<=818;
					out<=144;
				end
			end
			6685: begin
				if(in == 0) begin
					state<=6706;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=2817;
					out<=147;
				end
				if(in == 3) begin
					state<=4717;
					out<=148;
				end
				if(in == 4) begin
					state<=819;
					out<=149;
				end
			end
			6686: begin
				if(in == 0) begin
					state<=6697;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=2808;
					out<=152;
				end
				if(in == 3) begin
					state<=4708;
					out<=153;
				end
				if(in == 4) begin
					state<=810;
					out<=154;
				end
			end
			6687: begin
				if(in == 0) begin
					state<=7399;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=3510;
					out<=157;
				end
				if(in == 3) begin
					state<=5498;
					out<=158;
				end
				if(in == 4) begin
					state<=1609;
					out<=159;
				end
			end
			6688: begin
				if(in == 0) begin
					state<=7400;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=3511;
					out<=162;
				end
				if(in == 3) begin
					state<=5499;
					out<=163;
				end
				if(in == 4) begin
					state<=1610;
					out<=164;
				end
			end
			6689: begin
				if(in == 0) begin
					state<=7401;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=3512;
					out<=167;
				end
				if(in == 3) begin
					state<=5500;
					out<=168;
				end
				if(in == 4) begin
					state<=1611;
					out<=169;
				end
			end
			6690: begin
				if(in == 0) begin
					state<=7402;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=3513;
					out<=172;
				end
				if(in == 3) begin
					state<=5501;
					out<=173;
				end
				if(in == 4) begin
					state<=1612;
					out<=174;
				end
			end
			6691: begin
				if(in == 0) begin
					state<=7403;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=3514;
					out<=177;
				end
				if(in == 3) begin
					state<=5502;
					out<=178;
				end
				if(in == 4) begin
					state<=1613;
					out<=179;
				end
			end
			6692: begin
				if(in == 0) begin
					state<=7404;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=3515;
					out<=182;
				end
				if(in == 3) begin
					state<=5503;
					out<=183;
				end
				if(in == 4) begin
					state<=1614;
					out<=184;
				end
			end
			6693: begin
				if(in == 0) begin
					state<=7405;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=3516;
					out<=187;
				end
				if(in == 3) begin
					state<=5504;
					out<=188;
				end
				if(in == 4) begin
					state<=1615;
					out<=189;
				end
			end
			6694: begin
				if(in == 0) begin
					state<=7406;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=3517;
					out<=192;
				end
				if(in == 3) begin
					state<=5505;
					out<=193;
				end
				if(in == 4) begin
					state<=1616;
					out<=194;
				end
			end
			6695: begin
				if(in == 0) begin
					state<=7407;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=3518;
					out<=197;
				end
				if(in == 3) begin
					state<=5506;
					out<=198;
				end
				if(in == 4) begin
					state<=1617;
					out<=199;
				end
			end
			6696: begin
				if(in == 0) begin
					state<=7398;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=3509;
					out<=202;
				end
				if(in == 3) begin
					state<=5497;
					out<=203;
				end
				if(in == 4) begin
					state<=1608;
					out<=204;
				end
			end
			6697: begin
				if(in == 0) begin
					state<=6708;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=2819;
					out<=207;
				end
				if(in == 3) begin
					state<=4719;
					out<=208;
				end
				if(in == 4) begin
					state<=821;
					out<=209;
				end
			end
			6698: begin
				if(in == 0) begin
					state<=6709;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=2820;
					out<=212;
				end
				if(in == 3) begin
					state<=4720;
					out<=213;
				end
				if(in == 4) begin
					state<=822;
					out<=214;
				end
			end
			6699: begin
				if(in == 0) begin
					state<=6710;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=2821;
					out<=217;
				end
				if(in == 3) begin
					state<=4721;
					out<=218;
				end
				if(in == 4) begin
					state<=823;
					out<=219;
				end
			end
			6700: begin
				if(in == 0) begin
					state<=6711;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=2822;
					out<=222;
				end
				if(in == 3) begin
					state<=4722;
					out<=223;
				end
				if(in == 4) begin
					state<=824;
					out<=224;
				end
			end
			6701: begin
				if(in == 0) begin
					state<=6712;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=2823;
					out<=227;
				end
				if(in == 3) begin
					state<=4723;
					out<=228;
				end
				if(in == 4) begin
					state<=825;
					out<=229;
				end
			end
			6702: begin
				if(in == 0) begin
					state<=6713;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=2824;
					out<=232;
				end
				if(in == 3) begin
					state<=4724;
					out<=233;
				end
				if(in == 4) begin
					state<=826;
					out<=234;
				end
			end
			6703: begin
				if(in == 0) begin
					state<=6714;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=2825;
					out<=237;
				end
				if(in == 3) begin
					state<=4725;
					out<=238;
				end
				if(in == 4) begin
					state<=827;
					out<=239;
				end
			end
			6704: begin
				if(in == 0) begin
					state<=6715;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=2826;
					out<=242;
				end
				if(in == 3) begin
					state<=4726;
					out<=243;
				end
				if(in == 4) begin
					state<=828;
					out<=244;
				end
			end
			6705: begin
				if(in == 0) begin
					state<=6716;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=2827;
					out<=247;
				end
				if(in == 3) begin
					state<=4727;
					out<=248;
				end
				if(in == 4) begin
					state<=829;
					out<=249;
				end
			end
			6706: begin
				if(in == 0) begin
					state<=6707;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=2818;
					out<=252;
				end
				if(in == 3) begin
					state<=4718;
					out<=253;
				end
				if(in == 4) begin
					state<=820;
					out<=254;
				end
			end
			6707: begin
				if(in == 0) begin
					state<=6718;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=2829;
					out<=1;
				end
				if(in == 3) begin
					state<=4729;
					out<=2;
				end
				if(in == 4) begin
					state<=831;
					out<=3;
				end
			end
			6708: begin
				if(in == 0) begin
					state<=6719;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=2830;
					out<=6;
				end
				if(in == 3) begin
					state<=4730;
					out<=7;
				end
				if(in == 4) begin
					state<=832;
					out<=8;
				end
			end
			6709: begin
				if(in == 0) begin
					state<=6720;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=2831;
					out<=11;
				end
				if(in == 3) begin
					state<=4731;
					out<=12;
				end
				if(in == 4) begin
					state<=833;
					out<=13;
				end
			end
			6710: begin
				if(in == 0) begin
					state<=6721;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=2832;
					out<=16;
				end
				if(in == 3) begin
					state<=4732;
					out<=17;
				end
				if(in == 4) begin
					state<=834;
					out<=18;
				end
			end
			6711: begin
				if(in == 0) begin
					state<=6722;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=2833;
					out<=21;
				end
				if(in == 3) begin
					state<=4733;
					out<=22;
				end
				if(in == 4) begin
					state<=835;
					out<=23;
				end
			end
			6712: begin
				if(in == 0) begin
					state<=6723;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=2834;
					out<=26;
				end
				if(in == 3) begin
					state<=4734;
					out<=27;
				end
				if(in == 4) begin
					state<=836;
					out<=28;
				end
			end
			6713: begin
				if(in == 0) begin
					state<=6724;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=2835;
					out<=31;
				end
				if(in == 3) begin
					state<=4735;
					out<=32;
				end
				if(in == 4) begin
					state<=837;
					out<=33;
				end
			end
			6714: begin
				if(in == 0) begin
					state<=6725;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=2836;
					out<=36;
				end
				if(in == 3) begin
					state<=4736;
					out<=37;
				end
				if(in == 4) begin
					state<=838;
					out<=38;
				end
			end
			6715: begin
				if(in == 0) begin
					state<=6726;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=2837;
					out<=41;
				end
				if(in == 3) begin
					state<=4737;
					out<=42;
				end
				if(in == 4) begin
					state<=839;
					out<=43;
				end
			end
			6716: begin
				if(in == 0) begin
					state<=6717;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=2828;
					out<=46;
				end
				if(in == 3) begin
					state<=4728;
					out<=47;
				end
				if(in == 4) begin
					state<=830;
					out<=48;
				end
			end
			6717: begin
				if(in == 0) begin
					state<=6728;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=2839;
					out<=51;
				end
				if(in == 3) begin
					state<=4739;
					out<=52;
				end
				if(in == 4) begin
					state<=841;
					out<=53;
				end
			end
			6718: begin
				if(in == 0) begin
					state<=6729;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=2840;
					out<=56;
				end
				if(in == 3) begin
					state<=4740;
					out<=57;
				end
				if(in == 4) begin
					state<=842;
					out<=58;
				end
			end
			6719: begin
				if(in == 0) begin
					state<=6730;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=2841;
					out<=61;
				end
				if(in == 3) begin
					state<=4741;
					out<=62;
				end
				if(in == 4) begin
					state<=843;
					out<=63;
				end
			end
			6720: begin
				if(in == 0) begin
					state<=6731;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=2842;
					out<=66;
				end
				if(in == 3) begin
					state<=4742;
					out<=67;
				end
				if(in == 4) begin
					state<=844;
					out<=68;
				end
			end
			6721: begin
				if(in == 0) begin
					state<=6732;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=2843;
					out<=71;
				end
				if(in == 3) begin
					state<=4743;
					out<=72;
				end
				if(in == 4) begin
					state<=845;
					out<=73;
				end
			end
			6722: begin
				if(in == 0) begin
					state<=6733;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=2844;
					out<=76;
				end
				if(in == 3) begin
					state<=4744;
					out<=77;
				end
				if(in == 4) begin
					state<=846;
					out<=78;
				end
			end
			6723: begin
				if(in == 0) begin
					state<=6734;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=2845;
					out<=81;
				end
				if(in == 3) begin
					state<=4745;
					out<=82;
				end
				if(in == 4) begin
					state<=847;
					out<=83;
				end
			end
			6724: begin
				if(in == 0) begin
					state<=6735;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=2846;
					out<=86;
				end
				if(in == 3) begin
					state<=4746;
					out<=87;
				end
				if(in == 4) begin
					state<=848;
					out<=88;
				end
			end
			6725: begin
				if(in == 0) begin
					state<=6736;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=2847;
					out<=91;
				end
				if(in == 3) begin
					state<=4747;
					out<=92;
				end
				if(in == 4) begin
					state<=849;
					out<=93;
				end
			end
			6726: begin
				if(in == 0) begin
					state<=6727;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=2838;
					out<=96;
				end
				if(in == 3) begin
					state<=4738;
					out<=97;
				end
				if(in == 4) begin
					state<=840;
					out<=98;
				end
			end
			6727: begin
				if(in == 0) begin
					state<=6738;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=2849;
					out<=101;
				end
				if(in == 3) begin
					state<=4749;
					out<=102;
				end
				if(in == 4) begin
					state<=851;
					out<=103;
				end
			end
			6728: begin
				if(in == 0) begin
					state<=6739;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=2850;
					out<=106;
				end
				if(in == 3) begin
					state<=4750;
					out<=107;
				end
				if(in == 4) begin
					state<=852;
					out<=108;
				end
			end
			6729: begin
				if(in == 0) begin
					state<=6740;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=2851;
					out<=111;
				end
				if(in == 3) begin
					state<=4751;
					out<=112;
				end
				if(in == 4) begin
					state<=853;
					out<=113;
				end
			end
			6730: begin
				if(in == 0) begin
					state<=6741;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=2852;
					out<=116;
				end
				if(in == 3) begin
					state<=4752;
					out<=117;
				end
				if(in == 4) begin
					state<=854;
					out<=118;
				end
			end
			6731: begin
				if(in == 0) begin
					state<=6742;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=2853;
					out<=121;
				end
				if(in == 3) begin
					state<=4753;
					out<=122;
				end
				if(in == 4) begin
					state<=855;
					out<=123;
				end
			end
			6732: begin
				if(in == 0) begin
					state<=6743;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=2854;
					out<=126;
				end
				if(in == 3) begin
					state<=4754;
					out<=127;
				end
				if(in == 4) begin
					state<=856;
					out<=128;
				end
			end
			6733: begin
				if(in == 0) begin
					state<=6744;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=2855;
					out<=131;
				end
				if(in == 3) begin
					state<=4755;
					out<=132;
				end
				if(in == 4) begin
					state<=857;
					out<=133;
				end
			end
			6734: begin
				if(in == 0) begin
					state<=6745;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=2856;
					out<=136;
				end
				if(in == 3) begin
					state<=4756;
					out<=137;
				end
				if(in == 4) begin
					state<=858;
					out<=138;
				end
			end
			6735: begin
				if(in == 0) begin
					state<=6746;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=2857;
					out<=141;
				end
				if(in == 3) begin
					state<=4757;
					out<=142;
				end
				if(in == 4) begin
					state<=859;
					out<=143;
				end
			end
			6736: begin
				if(in == 0) begin
					state<=6737;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=2848;
					out<=146;
				end
				if(in == 3) begin
					state<=4748;
					out<=147;
				end
				if(in == 4) begin
					state<=850;
					out<=148;
				end
			end
			6737: begin
				if(in == 0) begin
					state<=6748;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=2859;
					out<=151;
				end
				if(in == 3) begin
					state<=4759;
					out<=152;
				end
				if(in == 4) begin
					state<=861;
					out<=153;
				end
			end
			6738: begin
				if(in == 0) begin
					state<=6749;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=2860;
					out<=156;
				end
				if(in == 3) begin
					state<=4760;
					out<=157;
				end
				if(in == 4) begin
					state<=862;
					out<=158;
				end
			end
			6739: begin
				if(in == 0) begin
					state<=6750;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=2861;
					out<=161;
				end
				if(in == 3) begin
					state<=4761;
					out<=162;
				end
				if(in == 4) begin
					state<=863;
					out<=163;
				end
			end
			6740: begin
				if(in == 0) begin
					state<=6751;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=2862;
					out<=166;
				end
				if(in == 3) begin
					state<=4762;
					out<=167;
				end
				if(in == 4) begin
					state<=864;
					out<=168;
				end
			end
			6741: begin
				if(in == 0) begin
					state<=6752;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=2863;
					out<=171;
				end
				if(in == 3) begin
					state<=4763;
					out<=172;
				end
				if(in == 4) begin
					state<=865;
					out<=173;
				end
			end
			6742: begin
				if(in == 0) begin
					state<=6753;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=2864;
					out<=176;
				end
				if(in == 3) begin
					state<=4764;
					out<=177;
				end
				if(in == 4) begin
					state<=866;
					out<=178;
				end
			end
			6743: begin
				if(in == 0) begin
					state<=6754;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=2865;
					out<=181;
				end
				if(in == 3) begin
					state<=4765;
					out<=182;
				end
				if(in == 4) begin
					state<=867;
					out<=183;
				end
			end
			6744: begin
				if(in == 0) begin
					state<=6755;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=2866;
					out<=186;
				end
				if(in == 3) begin
					state<=4766;
					out<=187;
				end
				if(in == 4) begin
					state<=868;
					out<=188;
				end
			end
			6745: begin
				if(in == 0) begin
					state<=6756;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=2867;
					out<=191;
				end
				if(in == 3) begin
					state<=4767;
					out<=192;
				end
				if(in == 4) begin
					state<=869;
					out<=193;
				end
			end
			6746: begin
				if(in == 0) begin
					state<=6747;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=2858;
					out<=196;
				end
				if(in == 3) begin
					state<=4758;
					out<=197;
				end
				if(in == 4) begin
					state<=860;
					out<=198;
				end
			end
			6747: begin
				if(in == 0) begin
					state<=6758;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=2869;
					out<=201;
				end
				if(in == 3) begin
					state<=4769;
					out<=202;
				end
				if(in == 4) begin
					state<=871;
					out<=203;
				end
			end
			6748: begin
				if(in == 0) begin
					state<=6759;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=2870;
					out<=206;
				end
				if(in == 3) begin
					state<=4770;
					out<=207;
				end
				if(in == 4) begin
					state<=872;
					out<=208;
				end
			end
			6749: begin
				if(in == 0) begin
					state<=6760;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=2871;
					out<=211;
				end
				if(in == 3) begin
					state<=4771;
					out<=212;
				end
				if(in == 4) begin
					state<=873;
					out<=213;
				end
			end
			6750: begin
				if(in == 0) begin
					state<=6761;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=2872;
					out<=216;
				end
				if(in == 3) begin
					state<=4772;
					out<=217;
				end
				if(in == 4) begin
					state<=874;
					out<=218;
				end
			end
			6751: begin
				if(in == 0) begin
					state<=6762;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=2873;
					out<=221;
				end
				if(in == 3) begin
					state<=4773;
					out<=222;
				end
				if(in == 4) begin
					state<=875;
					out<=223;
				end
			end
			6752: begin
				if(in == 0) begin
					state<=6763;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=2874;
					out<=226;
				end
				if(in == 3) begin
					state<=4774;
					out<=227;
				end
				if(in == 4) begin
					state<=876;
					out<=228;
				end
			end
			6753: begin
				if(in == 0) begin
					state<=6764;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=2875;
					out<=231;
				end
				if(in == 3) begin
					state<=4775;
					out<=232;
				end
				if(in == 4) begin
					state<=877;
					out<=233;
				end
			end
			6754: begin
				if(in == 0) begin
					state<=6765;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=2876;
					out<=236;
				end
				if(in == 3) begin
					state<=4776;
					out<=237;
				end
				if(in == 4) begin
					state<=878;
					out<=238;
				end
			end
			6755: begin
				if(in == 0) begin
					state<=6766;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=2877;
					out<=241;
				end
				if(in == 3) begin
					state<=4777;
					out<=242;
				end
				if(in == 4) begin
					state<=879;
					out<=243;
				end
			end
			6756: begin
				if(in == 0) begin
					state<=6757;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=2868;
					out<=246;
				end
				if(in == 3) begin
					state<=4768;
					out<=247;
				end
				if(in == 4) begin
					state<=870;
					out<=248;
				end
			end
			6757: begin
				if(in == 0) begin
					state<=6768;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=2879;
					out<=251;
				end
				if(in == 3) begin
					state<=4779;
					out<=252;
				end
				if(in == 4) begin
					state<=881;
					out<=253;
				end
			end
			6758: begin
				if(in == 0) begin
					state<=6769;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=2880;
					out<=0;
				end
				if(in == 3) begin
					state<=4780;
					out<=1;
				end
				if(in == 4) begin
					state<=882;
					out<=2;
				end
			end
			6759: begin
				if(in == 0) begin
					state<=6770;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=2881;
					out<=5;
				end
				if(in == 3) begin
					state<=4781;
					out<=6;
				end
				if(in == 4) begin
					state<=883;
					out<=7;
				end
			end
			6760: begin
				if(in == 0) begin
					state<=6771;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=2882;
					out<=10;
				end
				if(in == 3) begin
					state<=4782;
					out<=11;
				end
				if(in == 4) begin
					state<=884;
					out<=12;
				end
			end
			6761: begin
				if(in == 0) begin
					state<=6772;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=2883;
					out<=15;
				end
				if(in == 3) begin
					state<=4783;
					out<=16;
				end
				if(in == 4) begin
					state<=885;
					out<=17;
				end
			end
			6762: begin
				if(in == 0) begin
					state<=6773;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=2884;
					out<=20;
				end
				if(in == 3) begin
					state<=4784;
					out<=21;
				end
				if(in == 4) begin
					state<=886;
					out<=22;
				end
			end
			6763: begin
				if(in == 0) begin
					state<=6774;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=2885;
					out<=25;
				end
				if(in == 3) begin
					state<=4785;
					out<=26;
				end
				if(in == 4) begin
					state<=887;
					out<=27;
				end
			end
			6764: begin
				if(in == 0) begin
					state<=6775;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=2886;
					out<=30;
				end
				if(in == 3) begin
					state<=4786;
					out<=31;
				end
				if(in == 4) begin
					state<=888;
					out<=32;
				end
			end
			6765: begin
				if(in == 0) begin
					state<=6776;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=2887;
					out<=35;
				end
				if(in == 3) begin
					state<=4787;
					out<=36;
				end
				if(in == 4) begin
					state<=889;
					out<=37;
				end
			end
			6766: begin
				if(in == 0) begin
					state<=6767;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=2878;
					out<=40;
				end
				if(in == 3) begin
					state<=4778;
					out<=41;
				end
				if(in == 4) begin
					state<=880;
					out<=42;
				end
			end
			6767: begin
				if(in == 0) begin
					state<=6778;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=2889;
					out<=45;
				end
				if(in == 3) begin
					state<=4789;
					out<=46;
				end
				if(in == 4) begin
					state<=891;
					out<=47;
				end
			end
			6768: begin
				if(in == 0) begin
					state<=6779;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=2890;
					out<=50;
				end
				if(in == 3) begin
					state<=4790;
					out<=51;
				end
				if(in == 4) begin
					state<=892;
					out<=52;
				end
			end
			6769: begin
				if(in == 0) begin
					state<=6780;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=2891;
					out<=55;
				end
				if(in == 3) begin
					state<=4791;
					out<=56;
				end
				if(in == 4) begin
					state<=893;
					out<=57;
				end
			end
			6770: begin
				if(in == 0) begin
					state<=6781;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=2892;
					out<=60;
				end
				if(in == 3) begin
					state<=4792;
					out<=61;
				end
				if(in == 4) begin
					state<=894;
					out<=62;
				end
			end
			6771: begin
				if(in == 0) begin
					state<=6782;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=2893;
					out<=65;
				end
				if(in == 3) begin
					state<=4793;
					out<=66;
				end
				if(in == 4) begin
					state<=895;
					out<=67;
				end
			end
			6772: begin
				if(in == 0) begin
					state<=6783;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=2894;
					out<=70;
				end
				if(in == 3) begin
					state<=4794;
					out<=71;
				end
				if(in == 4) begin
					state<=896;
					out<=72;
				end
			end
			6773: begin
				if(in == 0) begin
					state<=6784;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=2895;
					out<=75;
				end
				if(in == 3) begin
					state<=4795;
					out<=76;
				end
				if(in == 4) begin
					state<=897;
					out<=77;
				end
			end
			6774: begin
				if(in == 0) begin
					state<=6785;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=2896;
					out<=80;
				end
				if(in == 3) begin
					state<=4796;
					out<=81;
				end
				if(in == 4) begin
					state<=898;
					out<=82;
				end
			end
			6775: begin
				if(in == 0) begin
					state<=6786;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=2897;
					out<=85;
				end
				if(in == 3) begin
					state<=4797;
					out<=86;
				end
				if(in == 4) begin
					state<=899;
					out<=87;
				end
			end
			6776: begin
				if(in == 0) begin
					state<=6777;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=2888;
					out<=90;
				end
				if(in == 3) begin
					state<=4788;
					out<=91;
				end
				if(in == 4) begin
					state<=890;
					out<=92;
				end
			end
			6777: begin
				if(in == 0) begin
					state<=6688;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=2799;
					out<=95;
				end
				if(in == 3) begin
					state<=4699;
					out<=96;
				end
				if(in == 4) begin
					state<=801;
					out<=97;
				end
			end
			6778: begin
				if(in == 0) begin
					state<=6689;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=2800;
					out<=100;
				end
				if(in == 3) begin
					state<=4700;
					out<=101;
				end
				if(in == 4) begin
					state<=802;
					out<=102;
				end
			end
			6779: begin
				if(in == 0) begin
					state<=6690;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=2801;
					out<=105;
				end
				if(in == 3) begin
					state<=4701;
					out<=106;
				end
				if(in == 4) begin
					state<=803;
					out<=107;
				end
			end
			6780: begin
				if(in == 0) begin
					state<=6691;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=2802;
					out<=110;
				end
				if(in == 3) begin
					state<=4702;
					out<=111;
				end
				if(in == 4) begin
					state<=804;
					out<=112;
				end
			end
			6781: begin
				if(in == 0) begin
					state<=6692;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=2803;
					out<=115;
				end
				if(in == 3) begin
					state<=4703;
					out<=116;
				end
				if(in == 4) begin
					state<=805;
					out<=117;
				end
			end
			6782: begin
				if(in == 0) begin
					state<=6693;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=2804;
					out<=120;
				end
				if(in == 3) begin
					state<=4704;
					out<=121;
				end
				if(in == 4) begin
					state<=806;
					out<=122;
				end
			end
			6783: begin
				if(in == 0) begin
					state<=6694;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=2805;
					out<=125;
				end
				if(in == 3) begin
					state<=4705;
					out<=126;
				end
				if(in == 4) begin
					state<=807;
					out<=127;
				end
			end
			6784: begin
				if(in == 0) begin
					state<=6695;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=2806;
					out<=130;
				end
				if(in == 3) begin
					state<=4706;
					out<=131;
				end
				if(in == 4) begin
					state<=808;
					out<=132;
				end
			end
			6785: begin
				if(in == 0) begin
					state<=6696;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=2807;
					out<=135;
				end
				if(in == 3) begin
					state<=4707;
					out<=136;
				end
				if(in == 4) begin
					state<=809;
					out<=137;
				end
			end
			6786: begin
				if(in == 0) begin
					state<=6687;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=2798;
					out<=140;
				end
				if(in == 3) begin
					state<=4698;
					out<=141;
				end
				if(in == 4) begin
					state<=800;
					out<=142;
				end
			end
			6787: begin
				if(in == 0) begin
					state<=6798;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=2909;
					out<=145;
				end
				if(in == 3) begin
					state<=5353;
					out<=146;
				end
				if(in == 4) begin
					state<=1464;
					out<=147;
				end
			end
			6788: begin
				if(in == 0) begin
					state<=6799;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=2910;
					out<=150;
				end
				if(in == 3) begin
					state<=5354;
					out<=151;
				end
				if(in == 4) begin
					state<=1465;
					out<=152;
				end
			end
			6789: begin
				if(in == 0) begin
					state<=6800;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=2911;
					out<=155;
				end
				if(in == 3) begin
					state<=5355;
					out<=156;
				end
				if(in == 4) begin
					state<=1466;
					out<=157;
				end
			end
			6790: begin
				if(in == 0) begin
					state<=6801;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=2912;
					out<=160;
				end
				if(in == 3) begin
					state<=5356;
					out<=161;
				end
				if(in == 4) begin
					state<=1467;
					out<=162;
				end
			end
			6791: begin
				if(in == 0) begin
					state<=6802;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=2913;
					out<=165;
				end
				if(in == 3) begin
					state<=5357;
					out<=166;
				end
				if(in == 4) begin
					state<=1468;
					out<=167;
				end
			end
			6792: begin
				if(in == 0) begin
					state<=6803;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=2914;
					out<=170;
				end
				if(in == 3) begin
					state<=5358;
					out<=171;
				end
				if(in == 4) begin
					state<=1469;
					out<=172;
				end
			end
			6793: begin
				if(in == 0) begin
					state<=6804;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=2915;
					out<=175;
				end
				if(in == 3) begin
					state<=5359;
					out<=176;
				end
				if(in == 4) begin
					state<=1470;
					out<=177;
				end
			end
			6794: begin
				if(in == 0) begin
					state<=6805;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=2916;
					out<=180;
				end
				if(in == 3) begin
					state<=5360;
					out<=181;
				end
				if(in == 4) begin
					state<=1471;
					out<=182;
				end
			end
			6795: begin
				if(in == 0) begin
					state<=6806;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=2917;
					out<=185;
				end
				if(in == 3) begin
					state<=5361;
					out<=186;
				end
				if(in == 4) begin
					state<=1472;
					out<=187;
				end
			end
			6796: begin
				if(in == 0) begin
					state<=6797;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=2908;
					out<=190;
				end
				if(in == 3) begin
					state<=5352;
					out<=191;
				end
				if(in == 4) begin
					state<=1463;
					out<=192;
				end
			end
			6797: begin
				if(in == 0) begin
					state<=6808;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=2919;
					out<=195;
				end
				if(in == 3) begin
					state<=5363;
					out<=196;
				end
				if(in == 4) begin
					state<=1474;
					out<=197;
				end
			end
			6798: begin
				if(in == 0) begin
					state<=6809;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=2920;
					out<=200;
				end
				if(in == 3) begin
					state<=5364;
					out<=201;
				end
				if(in == 4) begin
					state<=1475;
					out<=202;
				end
			end
			6799: begin
				if(in == 0) begin
					state<=6810;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=2921;
					out<=205;
				end
				if(in == 3) begin
					state<=5365;
					out<=206;
				end
				if(in == 4) begin
					state<=1476;
					out<=207;
				end
			end
			6800: begin
				if(in == 0) begin
					state<=6811;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=2922;
					out<=210;
				end
				if(in == 3) begin
					state<=5366;
					out<=211;
				end
				if(in == 4) begin
					state<=1477;
					out<=212;
				end
			end
			6801: begin
				if(in == 0) begin
					state<=6812;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=2923;
					out<=215;
				end
				if(in == 3) begin
					state<=5367;
					out<=216;
				end
				if(in == 4) begin
					state<=1478;
					out<=217;
				end
			end
			6802: begin
				if(in == 0) begin
					state<=6813;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=2924;
					out<=220;
				end
				if(in == 3) begin
					state<=5368;
					out<=221;
				end
				if(in == 4) begin
					state<=1479;
					out<=222;
				end
			end
			6803: begin
				if(in == 0) begin
					state<=6814;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=2925;
					out<=225;
				end
				if(in == 3) begin
					state<=5369;
					out<=226;
				end
				if(in == 4) begin
					state<=1480;
					out<=227;
				end
			end
			6804: begin
				if(in == 0) begin
					state<=6815;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=2926;
					out<=230;
				end
				if(in == 3) begin
					state<=5370;
					out<=231;
				end
				if(in == 4) begin
					state<=1481;
					out<=232;
				end
			end
			6805: begin
				if(in == 0) begin
					state<=6816;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=2927;
					out<=235;
				end
				if(in == 3) begin
					state<=5371;
					out<=236;
				end
				if(in == 4) begin
					state<=1482;
					out<=237;
				end
			end
			6806: begin
				if(in == 0) begin
					state<=6807;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=2918;
					out<=240;
				end
				if(in == 3) begin
					state<=5362;
					out<=241;
				end
				if(in == 4) begin
					state<=1473;
					out<=242;
				end
			end
			6807: begin
				if(in == 0) begin
					state<=6214;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=2325;
					out<=245;
				end
				if(in == 3) begin
					state<=4225;
					out<=246;
				end
				if(in == 4) begin
					state<=327;
					out<=247;
				end
			end
			6808: begin
				if(in == 0) begin
					state<=6215;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=2326;
					out<=250;
				end
				if(in == 3) begin
					state<=4226;
					out<=251;
				end
				if(in == 4) begin
					state<=328;
					out<=252;
				end
			end
			6809: begin
				if(in == 0) begin
					state<=6216;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=2327;
					out<=255;
				end
				if(in == 3) begin
					state<=4227;
					out<=0;
				end
				if(in == 4) begin
					state<=329;
					out<=1;
				end
			end
			6810: begin
				if(in == 0) begin
					state<=6217;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=2328;
					out<=4;
				end
				if(in == 3) begin
					state<=4228;
					out<=5;
				end
				if(in == 4) begin
					state<=330;
					out<=6;
				end
			end
			6811: begin
				if(in == 0) begin
					state<=6218;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=2329;
					out<=9;
				end
				if(in == 3) begin
					state<=4229;
					out<=10;
				end
				if(in == 4) begin
					state<=331;
					out<=11;
				end
			end
			6812: begin
				if(in == 0) begin
					state<=6219;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=2330;
					out<=14;
				end
				if(in == 3) begin
					state<=4230;
					out<=15;
				end
				if(in == 4) begin
					state<=332;
					out<=16;
				end
			end
			6813: begin
				if(in == 0) begin
					state<=6220;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=2331;
					out<=19;
				end
				if(in == 3) begin
					state<=4231;
					out<=20;
				end
				if(in == 4) begin
					state<=333;
					out<=21;
				end
			end
			6814: begin
				if(in == 0) begin
					state<=6221;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=2332;
					out<=24;
				end
				if(in == 3) begin
					state<=4232;
					out<=25;
				end
				if(in == 4) begin
					state<=334;
					out<=26;
				end
			end
			6815: begin
				if(in == 0) begin
					state<=6222;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=2333;
					out<=29;
				end
				if(in == 3) begin
					state<=4233;
					out<=30;
				end
				if(in == 4) begin
					state<=335;
					out<=31;
				end
			end
			6816: begin
				if(in == 0) begin
					state<=6817;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=2928;
					out<=34;
				end
				if(in == 3) begin
					state<=5372;
					out<=35;
				end
				if(in == 4) begin
					state<=1483;
					out<=36;
				end
			end
			6817: begin
				if(in == 0) begin
					state<=6224;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=2335;
					out<=39;
				end
				if(in == 3) begin
					state<=4235;
					out<=40;
				end
				if(in == 4) begin
					state<=337;
					out<=41;
				end
			end
			6818: begin
				if(in == 0) begin
					state<=6829;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=2940;
					out<=44;
				end
				if(in == 3) begin
					state<=4255;
					out<=45;
				end
				if(in == 4) begin
					state<=357;
					out<=46;
				end
			end
			6819: begin
				if(in == 0) begin
					state<=6830;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=2941;
					out<=49;
				end
				if(in == 3) begin
					state<=4256;
					out<=50;
				end
				if(in == 4) begin
					state<=358;
					out<=51;
				end
			end
			6820: begin
				if(in == 0) begin
					state<=6831;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=2942;
					out<=54;
				end
				if(in == 3) begin
					state<=4257;
					out<=55;
				end
				if(in == 4) begin
					state<=359;
					out<=56;
				end
			end
			6821: begin
				if(in == 0) begin
					state<=6832;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=2943;
					out<=59;
				end
				if(in == 3) begin
					state<=4258;
					out<=60;
				end
				if(in == 4) begin
					state<=360;
					out<=61;
				end
			end
			6822: begin
				if(in == 0) begin
					state<=6833;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=2944;
					out<=64;
				end
				if(in == 3) begin
					state<=4259;
					out<=65;
				end
				if(in == 4) begin
					state<=361;
					out<=66;
				end
			end
			6823: begin
				if(in == 0) begin
					state<=6834;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=2945;
					out<=69;
				end
				if(in == 3) begin
					state<=4260;
					out<=70;
				end
				if(in == 4) begin
					state<=362;
					out<=71;
				end
			end
			6824: begin
				if(in == 0) begin
					state<=6835;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=2946;
					out<=74;
				end
				if(in == 3) begin
					state<=4261;
					out<=75;
				end
				if(in == 4) begin
					state<=363;
					out<=76;
				end
			end
			6825: begin
				if(in == 0) begin
					state<=6836;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=2947;
					out<=79;
				end
				if(in == 3) begin
					state<=4262;
					out<=80;
				end
				if(in == 4) begin
					state<=364;
					out<=81;
				end
			end
			6826: begin
				if(in == 0) begin
					state<=6837;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=2948;
					out<=84;
				end
				if(in == 3) begin
					state<=4263;
					out<=85;
				end
				if(in == 4) begin
					state<=365;
					out<=86;
				end
			end
			6827: begin
				if(in == 0) begin
					state<=6828;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=2939;
					out<=89;
				end
				if(in == 3) begin
					state<=4254;
					out<=90;
				end
				if(in == 4) begin
					state<=356;
					out<=91;
				end
			end
			6828: begin
				if(in == 0) begin
					state<=6839;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=2950;
					out<=94;
				end
				if(in == 3) begin
					state<=4265;
					out<=95;
				end
				if(in == 4) begin
					state<=367;
					out<=96;
				end
			end
			6829: begin
				if(in == 0) begin
					state<=6840;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=2951;
					out<=99;
				end
				if(in == 3) begin
					state<=4266;
					out<=100;
				end
				if(in == 4) begin
					state<=368;
					out<=101;
				end
			end
			6830: begin
				if(in == 0) begin
					state<=6841;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=2952;
					out<=104;
				end
				if(in == 3) begin
					state<=4267;
					out<=105;
				end
				if(in == 4) begin
					state<=369;
					out<=106;
				end
			end
			6831: begin
				if(in == 0) begin
					state<=6842;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=2953;
					out<=109;
				end
				if(in == 3) begin
					state<=4268;
					out<=110;
				end
				if(in == 4) begin
					state<=370;
					out<=111;
				end
			end
			6832: begin
				if(in == 0) begin
					state<=6843;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=2954;
					out<=114;
				end
				if(in == 3) begin
					state<=4269;
					out<=115;
				end
				if(in == 4) begin
					state<=371;
					out<=116;
				end
			end
			6833: begin
				if(in == 0) begin
					state<=6844;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=2955;
					out<=119;
				end
				if(in == 3) begin
					state<=4270;
					out<=120;
				end
				if(in == 4) begin
					state<=372;
					out<=121;
				end
			end
			6834: begin
				if(in == 0) begin
					state<=6845;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=2956;
					out<=124;
				end
				if(in == 3) begin
					state<=4271;
					out<=125;
				end
				if(in == 4) begin
					state<=373;
					out<=126;
				end
			end
			6835: begin
				if(in == 0) begin
					state<=6846;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=2957;
					out<=129;
				end
				if(in == 3) begin
					state<=4272;
					out<=130;
				end
				if(in == 4) begin
					state<=374;
					out<=131;
				end
			end
			6836: begin
				if(in == 0) begin
					state<=6847;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=2958;
					out<=134;
				end
				if(in == 3) begin
					state<=4273;
					out<=135;
				end
				if(in == 4) begin
					state<=375;
					out<=136;
				end
			end
			6837: begin
				if(in == 0) begin
					state<=6838;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=2949;
					out<=139;
				end
				if(in == 3) begin
					state<=4264;
					out<=140;
				end
				if(in == 4) begin
					state<=366;
					out<=141;
				end
			end
			6838: begin
				if(in == 0) begin
					state<=6849;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=2960;
					out<=144;
				end
				if(in == 3) begin
					state<=4275;
					out<=145;
				end
				if(in == 4) begin
					state<=377;
					out<=146;
				end
			end
			6839: begin
				if(in == 0) begin
					state<=6850;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=2961;
					out<=149;
				end
				if(in == 3) begin
					state<=4276;
					out<=150;
				end
				if(in == 4) begin
					state<=378;
					out<=151;
				end
			end
			6840: begin
				if(in == 0) begin
					state<=6851;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=2962;
					out<=154;
				end
				if(in == 3) begin
					state<=4277;
					out<=155;
				end
				if(in == 4) begin
					state<=379;
					out<=156;
				end
			end
			6841: begin
				if(in == 0) begin
					state<=6852;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=2963;
					out<=159;
				end
				if(in == 3) begin
					state<=4278;
					out<=160;
				end
				if(in == 4) begin
					state<=380;
					out<=161;
				end
			end
			6842: begin
				if(in == 0) begin
					state<=6853;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=2964;
					out<=164;
				end
				if(in == 3) begin
					state<=4279;
					out<=165;
				end
				if(in == 4) begin
					state<=381;
					out<=166;
				end
			end
			6843: begin
				if(in == 0) begin
					state<=6854;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=2965;
					out<=169;
				end
				if(in == 3) begin
					state<=4280;
					out<=170;
				end
				if(in == 4) begin
					state<=382;
					out<=171;
				end
			end
			6844: begin
				if(in == 0) begin
					state<=6855;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=2966;
					out<=174;
				end
				if(in == 3) begin
					state<=4281;
					out<=175;
				end
				if(in == 4) begin
					state<=383;
					out<=176;
				end
			end
			6845: begin
				if(in == 0) begin
					state<=6856;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=2967;
					out<=179;
				end
				if(in == 3) begin
					state<=4282;
					out<=180;
				end
				if(in == 4) begin
					state<=384;
					out<=181;
				end
			end
			6846: begin
				if(in == 0) begin
					state<=6857;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=2968;
					out<=184;
				end
				if(in == 3) begin
					state<=4283;
					out<=185;
				end
				if(in == 4) begin
					state<=385;
					out<=186;
				end
			end
			6847: begin
				if(in == 0) begin
					state<=6848;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=2959;
					out<=189;
				end
				if(in == 3) begin
					state<=4274;
					out<=190;
				end
				if(in == 4) begin
					state<=376;
					out<=191;
				end
			end
			6848: begin
				if(in == 0) begin
					state<=6859;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=2970;
					out<=194;
				end
				if(in == 3) begin
					state<=4285;
					out<=195;
				end
				if(in == 4) begin
					state<=387;
					out<=196;
				end
			end
			6849: begin
				if(in == 0) begin
					state<=6860;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=2971;
					out<=199;
				end
				if(in == 3) begin
					state<=4286;
					out<=200;
				end
				if(in == 4) begin
					state<=388;
					out<=201;
				end
			end
			6850: begin
				if(in == 0) begin
					state<=6861;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=2972;
					out<=204;
				end
				if(in == 3) begin
					state<=4287;
					out<=205;
				end
				if(in == 4) begin
					state<=389;
					out<=206;
				end
			end
			6851: begin
				if(in == 0) begin
					state<=6862;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=2973;
					out<=209;
				end
				if(in == 3) begin
					state<=4288;
					out<=210;
				end
				if(in == 4) begin
					state<=390;
					out<=211;
				end
			end
			6852: begin
				if(in == 0) begin
					state<=6863;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=2974;
					out<=214;
				end
				if(in == 3) begin
					state<=4289;
					out<=215;
				end
				if(in == 4) begin
					state<=391;
					out<=216;
				end
			end
			6853: begin
				if(in == 0) begin
					state<=6864;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=2975;
					out<=219;
				end
				if(in == 3) begin
					state<=4290;
					out<=220;
				end
				if(in == 4) begin
					state<=392;
					out<=221;
				end
			end
			6854: begin
				if(in == 0) begin
					state<=6865;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=2976;
					out<=224;
				end
				if(in == 3) begin
					state<=4291;
					out<=225;
				end
				if(in == 4) begin
					state<=393;
					out<=226;
				end
			end
			6855: begin
				if(in == 0) begin
					state<=6866;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=2977;
					out<=229;
				end
				if(in == 3) begin
					state<=4292;
					out<=230;
				end
				if(in == 4) begin
					state<=394;
					out<=231;
				end
			end
			6856: begin
				if(in == 0) begin
					state<=6867;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=2978;
					out<=234;
				end
				if(in == 3) begin
					state<=4293;
					out<=235;
				end
				if(in == 4) begin
					state<=395;
					out<=236;
				end
			end
			6857: begin
				if(in == 0) begin
					state<=6858;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=2969;
					out<=239;
				end
				if(in == 3) begin
					state<=4284;
					out<=240;
				end
				if(in == 4) begin
					state<=386;
					out<=241;
				end
			end
			6858: begin
				if(in == 0) begin
					state<=6869;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=2980;
					out<=244;
				end
				if(in == 3) begin
					state<=4898;
					out<=245;
				end
				if(in == 4) begin
					state<=1000;
					out<=246;
				end
			end
			6859: begin
				if(in == 0) begin
					state<=6870;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=2981;
					out<=249;
				end
				if(in == 3) begin
					state<=4899;
					out<=250;
				end
				if(in == 4) begin
					state<=1001;
					out<=251;
				end
			end
			6860: begin
				if(in == 0) begin
					state<=6871;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=2982;
					out<=254;
				end
				if(in == 3) begin
					state<=4900;
					out<=255;
				end
				if(in == 4) begin
					state<=1002;
					out<=0;
				end
			end
			6861: begin
				if(in == 0) begin
					state<=6872;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=2983;
					out<=3;
				end
				if(in == 3) begin
					state<=4901;
					out<=4;
				end
				if(in == 4) begin
					state<=1003;
					out<=5;
				end
			end
			6862: begin
				if(in == 0) begin
					state<=6873;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=2984;
					out<=8;
				end
				if(in == 3) begin
					state<=4902;
					out<=9;
				end
				if(in == 4) begin
					state<=1004;
					out<=10;
				end
			end
			6863: begin
				if(in == 0) begin
					state<=6874;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=2985;
					out<=13;
				end
				if(in == 3) begin
					state<=4903;
					out<=14;
				end
				if(in == 4) begin
					state<=1005;
					out<=15;
				end
			end
			6864: begin
				if(in == 0) begin
					state<=6875;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=2986;
					out<=18;
				end
				if(in == 3) begin
					state<=4904;
					out<=19;
				end
				if(in == 4) begin
					state<=1006;
					out<=20;
				end
			end
			6865: begin
				if(in == 0) begin
					state<=6876;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=2987;
					out<=23;
				end
				if(in == 3) begin
					state<=4905;
					out<=24;
				end
				if(in == 4) begin
					state<=1007;
					out<=25;
				end
			end
			6866: begin
				if(in == 0) begin
					state<=6877;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=2988;
					out<=28;
				end
				if(in == 3) begin
					state<=4906;
					out<=29;
				end
				if(in == 4) begin
					state<=1008;
					out<=30;
				end
			end
			6867: begin
				if(in == 0) begin
					state<=6868;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=2979;
					out<=33;
				end
				if(in == 3) begin
					state<=4897;
					out<=34;
				end
				if(in == 4) begin
					state<=999;
					out<=35;
				end
			end
			6868: begin
				if(in == 0) begin
					state<=6879;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=2990;
					out<=38;
				end
				if(in == 3) begin
					state<=4908;
					out<=39;
				end
				if(in == 4) begin
					state<=1010;
					out<=40;
				end
			end
			6869: begin
				if(in == 0) begin
					state<=6880;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=2991;
					out<=43;
				end
				if(in == 3) begin
					state<=4909;
					out<=44;
				end
				if(in == 4) begin
					state<=1011;
					out<=45;
				end
			end
			6870: begin
				if(in == 0) begin
					state<=6881;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=2992;
					out<=48;
				end
				if(in == 3) begin
					state<=4910;
					out<=49;
				end
				if(in == 4) begin
					state<=1012;
					out<=50;
				end
			end
			6871: begin
				if(in == 0) begin
					state<=6882;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=2993;
					out<=53;
				end
				if(in == 3) begin
					state<=4911;
					out<=54;
				end
				if(in == 4) begin
					state<=1013;
					out<=55;
				end
			end
			6872: begin
				if(in == 0) begin
					state<=6883;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=2994;
					out<=58;
				end
				if(in == 3) begin
					state<=4912;
					out<=59;
				end
				if(in == 4) begin
					state<=1014;
					out<=60;
				end
			end
			6873: begin
				if(in == 0) begin
					state<=6884;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=2995;
					out<=63;
				end
				if(in == 3) begin
					state<=4913;
					out<=64;
				end
				if(in == 4) begin
					state<=1015;
					out<=65;
				end
			end
			6874: begin
				if(in == 0) begin
					state<=6885;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=2996;
					out<=68;
				end
				if(in == 3) begin
					state<=4914;
					out<=69;
				end
				if(in == 4) begin
					state<=1016;
					out<=70;
				end
			end
			6875: begin
				if(in == 0) begin
					state<=6886;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=2997;
					out<=73;
				end
				if(in == 3) begin
					state<=4915;
					out<=74;
				end
				if(in == 4) begin
					state<=1017;
					out<=75;
				end
			end
			6876: begin
				if(in == 0) begin
					state<=6887;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=2998;
					out<=78;
				end
				if(in == 3) begin
					state<=4916;
					out<=79;
				end
				if(in == 4) begin
					state<=1018;
					out<=80;
				end
			end
			6877: begin
				if(in == 0) begin
					state<=6878;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=2989;
					out<=83;
				end
				if(in == 3) begin
					state<=4907;
					out<=84;
				end
				if(in == 4) begin
					state<=1009;
					out<=85;
				end
			end
			6878: begin
				if(in == 0) begin
					state<=6889;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=3000;
					out<=88;
				end
				if(in == 3) begin
					state<=4918;
					out<=89;
				end
				if(in == 4) begin
					state<=1020;
					out<=90;
				end
			end
			6879: begin
				if(in == 0) begin
					state<=6890;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=3001;
					out<=93;
				end
				if(in == 3) begin
					state<=4919;
					out<=94;
				end
				if(in == 4) begin
					state<=1021;
					out<=95;
				end
			end
			6880: begin
				if(in == 0) begin
					state<=6891;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=3002;
					out<=98;
				end
				if(in == 3) begin
					state<=4920;
					out<=99;
				end
				if(in == 4) begin
					state<=1022;
					out<=100;
				end
			end
			6881: begin
				if(in == 0) begin
					state<=6892;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=3003;
					out<=103;
				end
				if(in == 3) begin
					state<=4921;
					out<=104;
				end
				if(in == 4) begin
					state<=1023;
					out<=105;
				end
			end
			6882: begin
				if(in == 0) begin
					state<=6893;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=3004;
					out<=108;
				end
				if(in == 3) begin
					state<=4922;
					out<=109;
				end
				if(in == 4) begin
					state<=1024;
					out<=110;
				end
			end
			6883: begin
				if(in == 0) begin
					state<=6894;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=3005;
					out<=113;
				end
				if(in == 3) begin
					state<=4923;
					out<=114;
				end
				if(in == 4) begin
					state<=1025;
					out<=115;
				end
			end
			6884: begin
				if(in == 0) begin
					state<=6895;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=3006;
					out<=118;
				end
				if(in == 3) begin
					state<=4924;
					out<=119;
				end
				if(in == 4) begin
					state<=1026;
					out<=120;
				end
			end
			6885: begin
				if(in == 0) begin
					state<=6896;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=3007;
					out<=123;
				end
				if(in == 3) begin
					state<=4925;
					out<=124;
				end
				if(in == 4) begin
					state<=1027;
					out<=125;
				end
			end
			6886: begin
				if(in == 0) begin
					state<=6897;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=3008;
					out<=128;
				end
				if(in == 3) begin
					state<=4926;
					out<=129;
				end
				if(in == 4) begin
					state<=1028;
					out<=130;
				end
			end
			6887: begin
				if(in == 0) begin
					state<=6888;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=2999;
					out<=133;
				end
				if(in == 3) begin
					state<=4917;
					out<=134;
				end
				if(in == 4) begin
					state<=1019;
					out<=135;
				end
			end
			6888: begin
				if(in == 0) begin
					state<=6899;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=3010;
					out<=138;
				end
				if(in == 3) begin
					state<=4294;
					out<=139;
				end
				if(in == 4) begin
					state<=396;
					out<=140;
				end
			end
			6889: begin
				if(in == 0) begin
					state<=6900;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=3011;
					out<=143;
				end
				if(in == 3) begin
					state<=4295;
					out<=144;
				end
				if(in == 4) begin
					state<=397;
					out<=145;
				end
			end
			6890: begin
				if(in == 0) begin
					state<=6901;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=3012;
					out<=148;
				end
				if(in == 3) begin
					state<=4296;
					out<=149;
				end
				if(in == 4) begin
					state<=398;
					out<=150;
				end
			end
			6891: begin
				if(in == 0) begin
					state<=6902;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=3013;
					out<=153;
				end
				if(in == 3) begin
					state<=4297;
					out<=154;
				end
				if(in == 4) begin
					state<=399;
					out<=155;
				end
			end
			6892: begin
				if(in == 0) begin
					state<=6903;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=3014;
					out<=158;
				end
				if(in == 3) begin
					state<=4298;
					out<=159;
				end
				if(in == 4) begin
					state<=400;
					out<=160;
				end
			end
			6893: begin
				if(in == 0) begin
					state<=6904;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=3015;
					out<=163;
				end
				if(in == 3) begin
					state<=4299;
					out<=164;
				end
				if(in == 4) begin
					state<=401;
					out<=165;
				end
			end
			6894: begin
				if(in == 0) begin
					state<=6905;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=3016;
					out<=168;
				end
				if(in == 3) begin
					state<=4300;
					out<=169;
				end
				if(in == 4) begin
					state<=402;
					out<=170;
				end
			end
			6895: begin
				if(in == 0) begin
					state<=6906;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=3017;
					out<=173;
				end
				if(in == 3) begin
					state<=4301;
					out<=174;
				end
				if(in == 4) begin
					state<=403;
					out<=175;
				end
			end
			6896: begin
				if(in == 0) begin
					state<=6907;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=3018;
					out<=178;
				end
				if(in == 3) begin
					state<=4302;
					out<=179;
				end
				if(in == 4) begin
					state<=404;
					out<=180;
				end
			end
			6897: begin
				if(in == 0) begin
					state<=6898;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=3009;
					out<=183;
				end
				if(in == 3) begin
					state<=4927;
					out<=184;
				end
				if(in == 4) begin
					state<=1029;
					out<=185;
				end
			end
			6898: begin
				if(in == 0) begin
					state<=6909;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=3020;
					out<=188;
				end
				if(in == 3) begin
					state<=4304;
					out<=189;
				end
				if(in == 4) begin
					state<=406;
					out<=190;
				end
			end
			6899: begin
				if(in == 0) begin
					state<=6910;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=3021;
					out<=193;
				end
				if(in == 3) begin
					state<=4305;
					out<=194;
				end
				if(in == 4) begin
					state<=407;
					out<=195;
				end
			end
			6900: begin
				if(in == 0) begin
					state<=6911;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=3022;
					out<=198;
				end
				if(in == 3) begin
					state<=4306;
					out<=199;
				end
				if(in == 4) begin
					state<=408;
					out<=200;
				end
			end
			6901: begin
				if(in == 0) begin
					state<=6912;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=3023;
					out<=203;
				end
				if(in == 3) begin
					state<=4307;
					out<=204;
				end
				if(in == 4) begin
					state<=409;
					out<=205;
				end
			end
			6902: begin
				if(in == 0) begin
					state<=6913;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=3024;
					out<=208;
				end
				if(in == 3) begin
					state<=4308;
					out<=209;
				end
				if(in == 4) begin
					state<=410;
					out<=210;
				end
			end
			6903: begin
				if(in == 0) begin
					state<=6914;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=3025;
					out<=213;
				end
				if(in == 3) begin
					state<=4309;
					out<=214;
				end
				if(in == 4) begin
					state<=411;
					out<=215;
				end
			end
			6904: begin
				if(in == 0) begin
					state<=6915;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=3026;
					out<=218;
				end
				if(in == 3) begin
					state<=4310;
					out<=219;
				end
				if(in == 4) begin
					state<=412;
					out<=220;
				end
			end
			6905: begin
				if(in == 0) begin
					state<=6916;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=3027;
					out<=223;
				end
				if(in == 3) begin
					state<=4311;
					out<=224;
				end
				if(in == 4) begin
					state<=413;
					out<=225;
				end
			end
			6906: begin
				if(in == 0) begin
					state<=6917;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=3028;
					out<=228;
				end
				if(in == 3) begin
					state<=4312;
					out<=229;
				end
				if(in == 4) begin
					state<=414;
					out<=230;
				end
			end
			6907: begin
				if(in == 0) begin
					state<=6908;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=3019;
					out<=233;
				end
				if(in == 3) begin
					state<=4303;
					out<=234;
				end
				if(in == 4) begin
					state<=405;
					out<=235;
				end
			end
			6908: begin
				if(in == 0) begin
					state<=6919;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=3030;
					out<=238;
				end
				if(in == 3) begin
					state<=4929;
					out<=239;
				end
				if(in == 4) begin
					state<=1031;
					out<=240;
				end
			end
			6909: begin
				if(in == 0) begin
					state<=6920;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=3031;
					out<=243;
				end
				if(in == 3) begin
					state<=4930;
					out<=244;
				end
				if(in == 4) begin
					state<=1032;
					out<=245;
				end
			end
			6910: begin
				if(in == 0) begin
					state<=6921;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=3032;
					out<=248;
				end
				if(in == 3) begin
					state<=4931;
					out<=249;
				end
				if(in == 4) begin
					state<=1033;
					out<=250;
				end
			end
			6911: begin
				if(in == 0) begin
					state<=6922;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=3033;
					out<=253;
				end
				if(in == 3) begin
					state<=4932;
					out<=254;
				end
				if(in == 4) begin
					state<=1034;
					out<=255;
				end
			end
			6912: begin
				if(in == 0) begin
					state<=6923;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=3034;
					out<=2;
				end
				if(in == 3) begin
					state<=4933;
					out<=3;
				end
				if(in == 4) begin
					state<=1035;
					out<=4;
				end
			end
			6913: begin
				if(in == 0) begin
					state<=6924;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=3035;
					out<=7;
				end
				if(in == 3) begin
					state<=4934;
					out<=8;
				end
				if(in == 4) begin
					state<=1036;
					out<=9;
				end
			end
			6914: begin
				if(in == 0) begin
					state<=6925;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=3036;
					out<=12;
				end
				if(in == 3) begin
					state<=4935;
					out<=13;
				end
				if(in == 4) begin
					state<=1037;
					out<=14;
				end
			end
			6915: begin
				if(in == 0) begin
					state<=6926;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=3037;
					out<=17;
				end
				if(in == 3) begin
					state<=4936;
					out<=18;
				end
				if(in == 4) begin
					state<=1038;
					out<=19;
				end
			end
			6916: begin
				if(in == 0) begin
					state<=6927;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=3038;
					out<=22;
				end
				if(in == 3) begin
					state<=4937;
					out<=23;
				end
				if(in == 4) begin
					state<=1039;
					out<=24;
				end
			end
			6917: begin
				if(in == 0) begin
					state<=6918;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=3029;
					out<=27;
				end
				if(in == 3) begin
					state<=4928;
					out<=28;
				end
				if(in == 4) begin
					state<=1030;
					out<=29;
				end
			end
			6918: begin
				if(in == 0) begin
					state<=6929;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=3040;
					out<=32;
				end
				if(in == 3) begin
					state<=4939;
					out<=33;
				end
				if(in == 4) begin
					state<=1041;
					out<=34;
				end
			end
			6919: begin
				if(in == 0) begin
					state<=6930;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=3041;
					out<=37;
				end
				if(in == 3) begin
					state<=4940;
					out<=38;
				end
				if(in == 4) begin
					state<=1042;
					out<=39;
				end
			end
			6920: begin
				if(in == 0) begin
					state<=6931;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=3042;
					out<=42;
				end
				if(in == 3) begin
					state<=4941;
					out<=43;
				end
				if(in == 4) begin
					state<=1043;
					out<=44;
				end
			end
			6921: begin
				if(in == 0) begin
					state<=6932;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=3043;
					out<=47;
				end
				if(in == 3) begin
					state<=4942;
					out<=48;
				end
				if(in == 4) begin
					state<=1044;
					out<=49;
				end
			end
			6922: begin
				if(in == 0) begin
					state<=6933;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=3044;
					out<=52;
				end
				if(in == 3) begin
					state<=4943;
					out<=53;
				end
				if(in == 4) begin
					state<=1045;
					out<=54;
				end
			end
			6923: begin
				if(in == 0) begin
					state<=6934;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=3045;
					out<=57;
				end
				if(in == 3) begin
					state<=4944;
					out<=58;
				end
				if(in == 4) begin
					state<=1046;
					out<=59;
				end
			end
			6924: begin
				if(in == 0) begin
					state<=6935;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=3046;
					out<=62;
				end
				if(in == 3) begin
					state<=4945;
					out<=63;
				end
				if(in == 4) begin
					state<=1047;
					out<=64;
				end
			end
			6925: begin
				if(in == 0) begin
					state<=6936;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=3047;
					out<=67;
				end
				if(in == 3) begin
					state<=4946;
					out<=68;
				end
				if(in == 4) begin
					state<=1048;
					out<=69;
				end
			end
			6926: begin
				if(in == 0) begin
					state<=6937;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=3048;
					out<=72;
				end
				if(in == 3) begin
					state<=4947;
					out<=73;
				end
				if(in == 4) begin
					state<=1049;
					out<=74;
				end
			end
			6927: begin
				if(in == 0) begin
					state<=6928;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=3039;
					out<=77;
				end
				if(in == 3) begin
					state<=4938;
					out<=78;
				end
				if(in == 4) begin
					state<=1040;
					out<=79;
				end
			end
			6928: begin
				if(in == 0) begin
					state<=6939;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=3050;
					out<=82;
				end
				if(in == 3) begin
					state<=4949;
					out<=83;
				end
				if(in == 4) begin
					state<=1051;
					out<=84;
				end
			end
			6929: begin
				if(in == 0) begin
					state<=6940;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=3051;
					out<=87;
				end
				if(in == 3) begin
					state<=4950;
					out<=88;
				end
				if(in == 4) begin
					state<=1052;
					out<=89;
				end
			end
			6930: begin
				if(in == 0) begin
					state<=6941;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=3052;
					out<=92;
				end
				if(in == 3) begin
					state<=4951;
					out<=93;
				end
				if(in == 4) begin
					state<=1053;
					out<=94;
				end
			end
			6931: begin
				if(in == 0) begin
					state<=6942;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=3053;
					out<=97;
				end
				if(in == 3) begin
					state<=4952;
					out<=98;
				end
				if(in == 4) begin
					state<=1054;
					out<=99;
				end
			end
			6932: begin
				if(in == 0) begin
					state<=6943;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=3054;
					out<=102;
				end
				if(in == 3) begin
					state<=4953;
					out<=103;
				end
				if(in == 4) begin
					state<=1055;
					out<=104;
				end
			end
			6933: begin
				if(in == 0) begin
					state<=6944;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=3055;
					out<=107;
				end
				if(in == 3) begin
					state<=4954;
					out<=108;
				end
				if(in == 4) begin
					state<=1056;
					out<=109;
				end
			end
			6934: begin
				if(in == 0) begin
					state<=6945;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=3056;
					out<=112;
				end
				if(in == 3) begin
					state<=4955;
					out<=113;
				end
				if(in == 4) begin
					state<=1057;
					out<=114;
				end
			end
			6935: begin
				if(in == 0) begin
					state<=6946;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=3057;
					out<=117;
				end
				if(in == 3) begin
					state<=4956;
					out<=118;
				end
				if(in == 4) begin
					state<=1058;
					out<=119;
				end
			end
			6936: begin
				if(in == 0) begin
					state<=6947;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=3058;
					out<=122;
				end
				if(in == 3) begin
					state<=4957;
					out<=123;
				end
				if(in == 4) begin
					state<=1059;
					out<=124;
				end
			end
			6937: begin
				if(in == 0) begin
					state<=6938;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=3049;
					out<=127;
				end
				if(in == 3) begin
					state<=4948;
					out<=128;
				end
				if(in == 4) begin
					state<=1050;
					out<=129;
				end
			end
			6938: begin
				if(in == 0) begin
					state<=6949;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=3060;
					out<=132;
				end
				if(in == 3) begin
					state<=4959;
					out<=133;
				end
				if(in == 4) begin
					state<=1061;
					out<=134;
				end
			end
			6939: begin
				if(in == 0) begin
					state<=6950;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=3061;
					out<=137;
				end
				if(in == 3) begin
					state<=4960;
					out<=138;
				end
				if(in == 4) begin
					state<=1062;
					out<=139;
				end
			end
			6940: begin
				if(in == 0) begin
					state<=6951;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=3062;
					out<=142;
				end
				if(in == 3) begin
					state<=4961;
					out<=143;
				end
				if(in == 4) begin
					state<=1063;
					out<=144;
				end
			end
			6941: begin
				if(in == 0) begin
					state<=6952;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=3063;
					out<=147;
				end
				if(in == 3) begin
					state<=4962;
					out<=148;
				end
				if(in == 4) begin
					state<=1064;
					out<=149;
				end
			end
			6942: begin
				if(in == 0) begin
					state<=6953;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=3064;
					out<=152;
				end
				if(in == 3) begin
					state<=4963;
					out<=153;
				end
				if(in == 4) begin
					state<=1065;
					out<=154;
				end
			end
			6943: begin
				if(in == 0) begin
					state<=6954;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=3065;
					out<=157;
				end
				if(in == 3) begin
					state<=4964;
					out<=158;
				end
				if(in == 4) begin
					state<=1066;
					out<=159;
				end
			end
			6944: begin
				if(in == 0) begin
					state<=6955;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=3066;
					out<=162;
				end
				if(in == 3) begin
					state<=4965;
					out<=163;
				end
				if(in == 4) begin
					state<=1067;
					out<=164;
				end
			end
			6945: begin
				if(in == 0) begin
					state<=6956;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=3067;
					out<=167;
				end
				if(in == 3) begin
					state<=4966;
					out<=168;
				end
				if(in == 4) begin
					state<=1068;
					out<=169;
				end
			end
			6946: begin
				if(in == 0) begin
					state<=6957;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=3068;
					out<=172;
				end
				if(in == 3) begin
					state<=4967;
					out<=173;
				end
				if(in == 4) begin
					state<=1069;
					out<=174;
				end
			end
			6947: begin
				if(in == 0) begin
					state<=6948;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=3059;
					out<=177;
				end
				if(in == 3) begin
					state<=4958;
					out<=178;
				end
				if(in == 4) begin
					state<=1060;
					out<=179;
				end
			end
			6948: begin
				if(in == 0) begin
					state<=6959;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=3070;
					out<=182;
				end
				if(in == 3) begin
					state<=4969;
					out<=183;
				end
				if(in == 4) begin
					state<=1071;
					out<=184;
				end
			end
			6949: begin
				if(in == 0) begin
					state<=6960;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=3071;
					out<=187;
				end
				if(in == 3) begin
					state<=4970;
					out<=188;
				end
				if(in == 4) begin
					state<=1072;
					out<=189;
				end
			end
			6950: begin
				if(in == 0) begin
					state<=6961;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=3072;
					out<=192;
				end
				if(in == 3) begin
					state<=4971;
					out<=193;
				end
				if(in == 4) begin
					state<=1073;
					out<=194;
				end
			end
			6951: begin
				if(in == 0) begin
					state<=6962;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=3073;
					out<=197;
				end
				if(in == 3) begin
					state<=4972;
					out<=198;
				end
				if(in == 4) begin
					state<=1074;
					out<=199;
				end
			end
			6952: begin
				if(in == 0) begin
					state<=6963;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=3074;
					out<=202;
				end
				if(in == 3) begin
					state<=4973;
					out<=203;
				end
				if(in == 4) begin
					state<=1075;
					out<=204;
				end
			end
			6953: begin
				if(in == 0) begin
					state<=6964;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=3075;
					out<=207;
				end
				if(in == 3) begin
					state<=4974;
					out<=208;
				end
				if(in == 4) begin
					state<=1076;
					out<=209;
				end
			end
			6954: begin
				if(in == 0) begin
					state<=6965;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=3076;
					out<=212;
				end
				if(in == 3) begin
					state<=4975;
					out<=213;
				end
				if(in == 4) begin
					state<=1077;
					out<=214;
				end
			end
			6955: begin
				if(in == 0) begin
					state<=6966;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=3077;
					out<=217;
				end
				if(in == 3) begin
					state<=4976;
					out<=218;
				end
				if(in == 4) begin
					state<=1078;
					out<=219;
				end
			end
			6956: begin
				if(in == 0) begin
					state<=6967;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=3078;
					out<=222;
				end
				if(in == 3) begin
					state<=4977;
					out<=223;
				end
				if(in == 4) begin
					state<=1079;
					out<=224;
				end
			end
			6957: begin
				if(in == 0) begin
					state<=6958;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=3069;
					out<=227;
				end
				if(in == 3) begin
					state<=4968;
					out<=228;
				end
				if(in == 4) begin
					state<=1070;
					out<=229;
				end
			end
			6958: begin
				if(in == 0) begin
					state<=6969;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=3080;
					out<=232;
				end
				if(in == 3) begin
					state<=4979;
					out<=233;
				end
				if(in == 4) begin
					state<=1081;
					out<=234;
				end
			end
			6959: begin
				if(in == 0) begin
					state<=6970;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=3081;
					out<=237;
				end
				if(in == 3) begin
					state<=4980;
					out<=238;
				end
				if(in == 4) begin
					state<=1082;
					out<=239;
				end
			end
			6960: begin
				if(in == 0) begin
					state<=6971;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=3082;
					out<=242;
				end
				if(in == 3) begin
					state<=4981;
					out<=243;
				end
				if(in == 4) begin
					state<=1083;
					out<=244;
				end
			end
			6961: begin
				if(in == 0) begin
					state<=6972;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=3083;
					out<=247;
				end
				if(in == 3) begin
					state<=4982;
					out<=248;
				end
				if(in == 4) begin
					state<=1084;
					out<=249;
				end
			end
			6962: begin
				if(in == 0) begin
					state<=6973;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=3084;
					out<=252;
				end
				if(in == 3) begin
					state<=4983;
					out<=253;
				end
				if(in == 4) begin
					state<=1085;
					out<=254;
				end
			end
			6963: begin
				if(in == 0) begin
					state<=6974;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=3085;
					out<=1;
				end
				if(in == 3) begin
					state<=4984;
					out<=2;
				end
				if(in == 4) begin
					state<=1086;
					out<=3;
				end
			end
			6964: begin
				if(in == 0) begin
					state<=6975;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=3086;
					out<=6;
				end
				if(in == 3) begin
					state<=4985;
					out<=7;
				end
				if(in == 4) begin
					state<=1087;
					out<=8;
				end
			end
			6965: begin
				if(in == 0) begin
					state<=6976;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=3087;
					out<=11;
				end
				if(in == 3) begin
					state<=4986;
					out<=12;
				end
				if(in == 4) begin
					state<=1088;
					out<=13;
				end
			end
			6966: begin
				if(in == 0) begin
					state<=6977;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=3088;
					out<=16;
				end
				if(in == 3) begin
					state<=4987;
					out<=17;
				end
				if(in == 4) begin
					state<=1089;
					out<=18;
				end
			end
			6967: begin
				if(in == 0) begin
					state<=6968;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=3079;
					out<=21;
				end
				if(in == 3) begin
					state<=4978;
					out<=22;
				end
				if(in == 4) begin
					state<=1080;
					out<=23;
				end
			end
			6968: begin
				if(in == 0) begin
					state<=6979;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=3090;
					out<=26;
				end
				if(in == 3) begin
					state<=4989;
					out<=27;
				end
				if(in == 4) begin
					state<=1091;
					out<=28;
				end
			end
			6969: begin
				if(in == 0) begin
					state<=6980;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=3091;
					out<=31;
				end
				if(in == 3) begin
					state<=4990;
					out<=32;
				end
				if(in == 4) begin
					state<=1092;
					out<=33;
				end
			end
			6970: begin
				if(in == 0) begin
					state<=6981;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=3092;
					out<=36;
				end
				if(in == 3) begin
					state<=4991;
					out<=37;
				end
				if(in == 4) begin
					state<=1093;
					out<=38;
				end
			end
			6971: begin
				if(in == 0) begin
					state<=6982;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=3093;
					out<=41;
				end
				if(in == 3) begin
					state<=4992;
					out<=42;
				end
				if(in == 4) begin
					state<=1094;
					out<=43;
				end
			end
			6972: begin
				if(in == 0) begin
					state<=6983;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=3094;
					out<=46;
				end
				if(in == 3) begin
					state<=4993;
					out<=47;
				end
				if(in == 4) begin
					state<=1095;
					out<=48;
				end
			end
			6973: begin
				if(in == 0) begin
					state<=6984;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=3095;
					out<=51;
				end
				if(in == 3) begin
					state<=4994;
					out<=52;
				end
				if(in == 4) begin
					state<=1096;
					out<=53;
				end
			end
			6974: begin
				if(in == 0) begin
					state<=6985;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=3096;
					out<=56;
				end
				if(in == 3) begin
					state<=4995;
					out<=57;
				end
				if(in == 4) begin
					state<=1097;
					out<=58;
				end
			end
			6975: begin
				if(in == 0) begin
					state<=6986;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=3097;
					out<=61;
				end
				if(in == 3) begin
					state<=4996;
					out<=62;
				end
				if(in == 4) begin
					state<=1098;
					out<=63;
				end
			end
			6976: begin
				if(in == 0) begin
					state<=6987;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=3098;
					out<=66;
				end
				if(in == 3) begin
					state<=4997;
					out<=67;
				end
				if(in == 4) begin
					state<=1099;
					out<=68;
				end
			end
			6977: begin
				if(in == 0) begin
					state<=6978;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=3089;
					out<=71;
				end
				if(in == 3) begin
					state<=4988;
					out<=72;
				end
				if(in == 4) begin
					state<=1090;
					out<=73;
				end
			end
			6978: begin
				if(in == 0) begin
					state<=6989;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=3100;
					out<=76;
				end
				if(in == 3) begin
					state<=4999;
					out<=77;
				end
				if(in == 4) begin
					state<=1101;
					out<=78;
				end
			end
			6979: begin
				if(in == 0) begin
					state<=6990;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=3101;
					out<=81;
				end
				if(in == 3) begin
					state<=5000;
					out<=82;
				end
				if(in == 4) begin
					state<=1102;
					out<=83;
				end
			end
			6980: begin
				if(in == 0) begin
					state<=6991;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=3102;
					out<=86;
				end
				if(in == 3) begin
					state<=5001;
					out<=87;
				end
				if(in == 4) begin
					state<=1103;
					out<=88;
				end
			end
			6981: begin
				if(in == 0) begin
					state<=6992;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=3103;
					out<=91;
				end
				if(in == 3) begin
					state<=5002;
					out<=92;
				end
				if(in == 4) begin
					state<=1104;
					out<=93;
				end
			end
			6982: begin
				if(in == 0) begin
					state<=6993;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=3104;
					out<=96;
				end
				if(in == 3) begin
					state<=5003;
					out<=97;
				end
				if(in == 4) begin
					state<=1105;
					out<=98;
				end
			end
			6983: begin
				if(in == 0) begin
					state<=6994;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=3105;
					out<=101;
				end
				if(in == 3) begin
					state<=5004;
					out<=102;
				end
				if(in == 4) begin
					state<=1106;
					out<=103;
				end
			end
			6984: begin
				if(in == 0) begin
					state<=6995;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=3106;
					out<=106;
				end
				if(in == 3) begin
					state<=5005;
					out<=107;
				end
				if(in == 4) begin
					state<=1107;
					out<=108;
				end
			end
			6985: begin
				if(in == 0) begin
					state<=6996;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=3107;
					out<=111;
				end
				if(in == 3) begin
					state<=5006;
					out<=112;
				end
				if(in == 4) begin
					state<=1108;
					out<=113;
				end
			end
			6986: begin
				if(in == 0) begin
					state<=6997;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=3108;
					out<=116;
				end
				if(in == 3) begin
					state<=5007;
					out<=117;
				end
				if(in == 4) begin
					state<=1109;
					out<=118;
				end
			end
			6987: begin
				if(in == 0) begin
					state<=6988;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=3099;
					out<=121;
				end
				if(in == 3) begin
					state<=4998;
					out<=122;
				end
				if(in == 4) begin
					state<=1100;
					out<=123;
				end
			end
			6988: begin
				if(in == 0) begin
					state<=6999;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=3110;
					out<=126;
				end
				if(in == 3) begin
					state<=5009;
					out<=127;
				end
				if(in == 4) begin
					state<=1111;
					out<=128;
				end
			end
			6989: begin
				if(in == 0) begin
					state<=7000;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=3111;
					out<=131;
				end
				if(in == 3) begin
					state<=5010;
					out<=132;
				end
				if(in == 4) begin
					state<=1112;
					out<=133;
				end
			end
			6990: begin
				if(in == 0) begin
					state<=7001;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=3112;
					out<=136;
				end
				if(in == 3) begin
					state<=5011;
					out<=137;
				end
				if(in == 4) begin
					state<=1113;
					out<=138;
				end
			end
			6991: begin
				if(in == 0) begin
					state<=7002;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=3113;
					out<=141;
				end
				if(in == 3) begin
					state<=5012;
					out<=142;
				end
				if(in == 4) begin
					state<=1114;
					out<=143;
				end
			end
			6992: begin
				if(in == 0) begin
					state<=7003;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=3114;
					out<=146;
				end
				if(in == 3) begin
					state<=5013;
					out<=147;
				end
				if(in == 4) begin
					state<=1115;
					out<=148;
				end
			end
			6993: begin
				if(in == 0) begin
					state<=7004;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=3115;
					out<=151;
				end
				if(in == 3) begin
					state<=5014;
					out<=152;
				end
				if(in == 4) begin
					state<=1116;
					out<=153;
				end
			end
			6994: begin
				if(in == 0) begin
					state<=7005;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=3116;
					out<=156;
				end
				if(in == 3) begin
					state<=5015;
					out<=157;
				end
				if(in == 4) begin
					state<=1117;
					out<=158;
				end
			end
			6995: begin
				if(in == 0) begin
					state<=7006;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=3117;
					out<=161;
				end
				if(in == 3) begin
					state<=5016;
					out<=162;
				end
				if(in == 4) begin
					state<=1118;
					out<=163;
				end
			end
			6996: begin
				if(in == 0) begin
					state<=7007;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=3118;
					out<=166;
				end
				if(in == 3) begin
					state<=5017;
					out<=167;
				end
				if(in == 4) begin
					state<=1119;
					out<=168;
				end
			end
			6997: begin
				if(in == 0) begin
					state<=6998;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=3109;
					out<=171;
				end
				if(in == 3) begin
					state<=5008;
					out<=172;
				end
				if(in == 4) begin
					state<=1110;
					out<=173;
				end
			end
			6998: begin
				if(in == 0) begin
					state<=7009;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=3120;
					out<=176;
				end
				if(in == 3) begin
					state<=5019;
					out<=177;
				end
				if(in == 4) begin
					state<=1121;
					out<=178;
				end
			end
			6999: begin
				if(in == 0) begin
					state<=7010;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=3121;
					out<=181;
				end
				if(in == 3) begin
					state<=5020;
					out<=182;
				end
				if(in == 4) begin
					state<=1122;
					out<=183;
				end
			end
			7000: begin
				if(in == 0) begin
					state<=7011;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=3122;
					out<=186;
				end
				if(in == 3) begin
					state<=5021;
					out<=187;
				end
				if(in == 4) begin
					state<=1123;
					out<=188;
				end
			end
			7001: begin
				if(in == 0) begin
					state<=7012;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=3123;
					out<=191;
				end
				if(in == 3) begin
					state<=5022;
					out<=192;
				end
				if(in == 4) begin
					state<=1124;
					out<=193;
				end
			end
			7002: begin
				if(in == 0) begin
					state<=7013;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=3124;
					out<=196;
				end
				if(in == 3) begin
					state<=5023;
					out<=197;
				end
				if(in == 4) begin
					state<=1125;
					out<=198;
				end
			end
			7003: begin
				if(in == 0) begin
					state<=7014;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=3125;
					out<=201;
				end
				if(in == 3) begin
					state<=5024;
					out<=202;
				end
				if(in == 4) begin
					state<=1126;
					out<=203;
				end
			end
			7004: begin
				if(in == 0) begin
					state<=7015;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=3126;
					out<=206;
				end
				if(in == 3) begin
					state<=5025;
					out<=207;
				end
				if(in == 4) begin
					state<=1127;
					out<=208;
				end
			end
			7005: begin
				if(in == 0) begin
					state<=7016;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=3127;
					out<=211;
				end
				if(in == 3) begin
					state<=5026;
					out<=212;
				end
				if(in == 4) begin
					state<=1128;
					out<=213;
				end
			end
			7006: begin
				if(in == 0) begin
					state<=7017;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=3128;
					out<=216;
				end
				if(in == 3) begin
					state<=5027;
					out<=217;
				end
				if(in == 4) begin
					state<=1129;
					out<=218;
				end
			end
			7007: begin
				if(in == 0) begin
					state<=7008;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=3119;
					out<=221;
				end
				if(in == 3) begin
					state<=5018;
					out<=222;
				end
				if(in == 4) begin
					state<=1120;
					out<=223;
				end
			end
			7008: begin
				if(in == 0) begin
					state<=7019;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=3130;
					out<=226;
				end
				if(in == 3) begin
					state<=5029;
					out<=227;
				end
				if(in == 4) begin
					state<=1131;
					out<=228;
				end
			end
			7009: begin
				if(in == 0) begin
					state<=7020;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=3131;
					out<=231;
				end
				if(in == 3) begin
					state<=5030;
					out<=232;
				end
				if(in == 4) begin
					state<=1132;
					out<=233;
				end
			end
			7010: begin
				if(in == 0) begin
					state<=7021;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=3132;
					out<=236;
				end
				if(in == 3) begin
					state<=5031;
					out<=237;
				end
				if(in == 4) begin
					state<=1133;
					out<=238;
				end
			end
			7011: begin
				if(in == 0) begin
					state<=7022;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=3133;
					out<=241;
				end
				if(in == 3) begin
					state<=5032;
					out<=242;
				end
				if(in == 4) begin
					state<=1134;
					out<=243;
				end
			end
			7012: begin
				if(in == 0) begin
					state<=7023;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=3134;
					out<=246;
				end
				if(in == 3) begin
					state<=5033;
					out<=247;
				end
				if(in == 4) begin
					state<=1135;
					out<=248;
				end
			end
			7013: begin
				if(in == 0) begin
					state<=7024;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=3135;
					out<=251;
				end
				if(in == 3) begin
					state<=5034;
					out<=252;
				end
				if(in == 4) begin
					state<=1136;
					out<=253;
				end
			end
			7014: begin
				if(in == 0) begin
					state<=7025;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=3136;
					out<=0;
				end
				if(in == 3) begin
					state<=5035;
					out<=1;
				end
				if(in == 4) begin
					state<=1137;
					out<=2;
				end
			end
			7015: begin
				if(in == 0) begin
					state<=7026;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=3137;
					out<=5;
				end
				if(in == 3) begin
					state<=5036;
					out<=6;
				end
				if(in == 4) begin
					state<=1138;
					out<=7;
				end
			end
			7016: begin
				if(in == 0) begin
					state<=7027;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=3138;
					out<=10;
				end
				if(in == 3) begin
					state<=5037;
					out<=11;
				end
				if(in == 4) begin
					state<=1139;
					out<=12;
				end
			end
			7017: begin
				if(in == 0) begin
					state<=7018;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=3129;
					out<=15;
				end
				if(in == 3) begin
					state<=5028;
					out<=16;
				end
				if(in == 4) begin
					state<=1130;
					out<=17;
				end
			end
			7018: begin
				if(in == 0) begin
					state<=7029;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=3140;
					out<=20;
				end
				if(in == 3) begin
					state<=5039;
					out<=21;
				end
				if(in == 4) begin
					state<=1141;
					out<=22;
				end
			end
			7019: begin
				if(in == 0) begin
					state<=7030;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=3141;
					out<=25;
				end
				if(in == 3) begin
					state<=5040;
					out<=26;
				end
				if(in == 4) begin
					state<=1142;
					out<=27;
				end
			end
			7020: begin
				if(in == 0) begin
					state<=7031;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=3142;
					out<=30;
				end
				if(in == 3) begin
					state<=5041;
					out<=31;
				end
				if(in == 4) begin
					state<=1143;
					out<=32;
				end
			end
			7021: begin
				if(in == 0) begin
					state<=7032;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=3143;
					out<=35;
				end
				if(in == 3) begin
					state<=5042;
					out<=36;
				end
				if(in == 4) begin
					state<=1144;
					out<=37;
				end
			end
			7022: begin
				if(in == 0) begin
					state<=7033;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=3144;
					out<=40;
				end
				if(in == 3) begin
					state<=5043;
					out<=41;
				end
				if(in == 4) begin
					state<=1145;
					out<=42;
				end
			end
			7023: begin
				if(in == 0) begin
					state<=7034;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=3145;
					out<=45;
				end
				if(in == 3) begin
					state<=5044;
					out<=46;
				end
				if(in == 4) begin
					state<=1146;
					out<=47;
				end
			end
			7024: begin
				if(in == 0) begin
					state<=7035;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=3146;
					out<=50;
				end
				if(in == 3) begin
					state<=5045;
					out<=51;
				end
				if(in == 4) begin
					state<=1147;
					out<=52;
				end
			end
			7025: begin
				if(in == 0) begin
					state<=7036;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=3147;
					out<=55;
				end
				if(in == 3) begin
					state<=5046;
					out<=56;
				end
				if(in == 4) begin
					state<=1148;
					out<=57;
				end
			end
			7026: begin
				if(in == 0) begin
					state<=7037;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=3148;
					out<=60;
				end
				if(in == 3) begin
					state<=5047;
					out<=61;
				end
				if(in == 4) begin
					state<=1149;
					out<=62;
				end
			end
			7027: begin
				if(in == 0) begin
					state<=7028;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=3139;
					out<=65;
				end
				if(in == 3) begin
					state<=5038;
					out<=66;
				end
				if(in == 4) begin
					state<=1140;
					out<=67;
				end
			end
			7028: begin
				if(in == 0) begin
					state<=7039;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=3150;
					out<=70;
				end
				if(in == 3) begin
					state<=5049;
					out<=71;
				end
				if(in == 4) begin
					state<=1151;
					out<=72;
				end
			end
			7029: begin
				if(in == 0) begin
					state<=7040;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=3151;
					out<=75;
				end
				if(in == 3) begin
					state<=5050;
					out<=76;
				end
				if(in == 4) begin
					state<=1152;
					out<=77;
				end
			end
			7030: begin
				if(in == 0) begin
					state<=7041;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=3152;
					out<=80;
				end
				if(in == 3) begin
					state<=5051;
					out<=81;
				end
				if(in == 4) begin
					state<=1153;
					out<=82;
				end
			end
			7031: begin
				if(in == 0) begin
					state<=7042;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=3153;
					out<=85;
				end
				if(in == 3) begin
					state<=5052;
					out<=86;
				end
				if(in == 4) begin
					state<=1154;
					out<=87;
				end
			end
			7032: begin
				if(in == 0) begin
					state<=7043;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=3154;
					out<=90;
				end
				if(in == 3) begin
					state<=5053;
					out<=91;
				end
				if(in == 4) begin
					state<=1155;
					out<=92;
				end
			end
			7033: begin
				if(in == 0) begin
					state<=7044;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=3155;
					out<=95;
				end
				if(in == 3) begin
					state<=5054;
					out<=96;
				end
				if(in == 4) begin
					state<=1156;
					out<=97;
				end
			end
			7034: begin
				if(in == 0) begin
					state<=7045;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=3156;
					out<=100;
				end
				if(in == 3) begin
					state<=5055;
					out<=101;
				end
				if(in == 4) begin
					state<=1157;
					out<=102;
				end
			end
			7035: begin
				if(in == 0) begin
					state<=7046;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=3157;
					out<=105;
				end
				if(in == 3) begin
					state<=5056;
					out<=106;
				end
				if(in == 4) begin
					state<=1158;
					out<=107;
				end
			end
			7036: begin
				if(in == 0) begin
					state<=7047;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=3158;
					out<=110;
				end
				if(in == 3) begin
					state<=5057;
					out<=111;
				end
				if(in == 4) begin
					state<=1159;
					out<=112;
				end
			end
			7037: begin
				if(in == 0) begin
					state<=7038;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=3149;
					out<=115;
				end
				if(in == 3) begin
					state<=5048;
					out<=116;
				end
				if(in == 4) begin
					state<=1150;
					out<=117;
				end
			end
			7038: begin
				if(in == 0) begin
					state<=7049;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=3160;
					out<=120;
				end
				if(in == 3) begin
					state<=5059;
					out<=121;
				end
				if(in == 4) begin
					state<=1161;
					out<=122;
				end
			end
			7039: begin
				if(in == 0) begin
					state<=7050;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=3161;
					out<=125;
				end
				if(in == 3) begin
					state<=5060;
					out<=126;
				end
				if(in == 4) begin
					state<=1162;
					out<=127;
				end
			end
			7040: begin
				if(in == 0) begin
					state<=7051;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=3162;
					out<=130;
				end
				if(in == 3) begin
					state<=5061;
					out<=131;
				end
				if(in == 4) begin
					state<=1163;
					out<=132;
				end
			end
			7041: begin
				if(in == 0) begin
					state<=7052;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=3163;
					out<=135;
				end
				if(in == 3) begin
					state<=5062;
					out<=136;
				end
				if(in == 4) begin
					state<=1164;
					out<=137;
				end
			end
			7042: begin
				if(in == 0) begin
					state<=7053;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=3164;
					out<=140;
				end
				if(in == 3) begin
					state<=5063;
					out<=141;
				end
				if(in == 4) begin
					state<=1165;
					out<=142;
				end
			end
			7043: begin
				if(in == 0) begin
					state<=7054;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=3165;
					out<=145;
				end
				if(in == 3) begin
					state<=5064;
					out<=146;
				end
				if(in == 4) begin
					state<=1166;
					out<=147;
				end
			end
			7044: begin
				if(in == 0) begin
					state<=7055;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=3166;
					out<=150;
				end
				if(in == 3) begin
					state<=5065;
					out<=151;
				end
				if(in == 4) begin
					state<=1167;
					out<=152;
				end
			end
			7045: begin
				if(in == 0) begin
					state<=7056;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=3167;
					out<=155;
				end
				if(in == 3) begin
					state<=5066;
					out<=156;
				end
				if(in == 4) begin
					state<=1168;
					out<=157;
				end
			end
			7046: begin
				if(in == 0) begin
					state<=7057;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=3168;
					out<=160;
				end
				if(in == 3) begin
					state<=5067;
					out<=161;
				end
				if(in == 4) begin
					state<=1169;
					out<=162;
				end
			end
			7047: begin
				if(in == 0) begin
					state<=7048;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=3159;
					out<=165;
				end
				if(in == 3) begin
					state<=5058;
					out<=166;
				end
				if(in == 4) begin
					state<=1160;
					out<=167;
				end
			end
			7048: begin
				if(in == 0) begin
					state<=7059;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=3170;
					out<=170;
				end
				if(in == 3) begin
					state<=5069;
					out<=171;
				end
				if(in == 4) begin
					state<=1171;
					out<=172;
				end
			end
			7049: begin
				if(in == 0) begin
					state<=7060;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=3171;
					out<=175;
				end
				if(in == 3) begin
					state<=5070;
					out<=176;
				end
				if(in == 4) begin
					state<=1172;
					out<=177;
				end
			end
			7050: begin
				if(in == 0) begin
					state<=7061;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=3172;
					out<=180;
				end
				if(in == 3) begin
					state<=5071;
					out<=181;
				end
				if(in == 4) begin
					state<=1173;
					out<=182;
				end
			end
			7051: begin
				if(in == 0) begin
					state<=7062;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=3173;
					out<=185;
				end
				if(in == 3) begin
					state<=5072;
					out<=186;
				end
				if(in == 4) begin
					state<=1174;
					out<=187;
				end
			end
			7052: begin
				if(in == 0) begin
					state<=7063;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=3174;
					out<=190;
				end
				if(in == 3) begin
					state<=5073;
					out<=191;
				end
				if(in == 4) begin
					state<=1175;
					out<=192;
				end
			end
			7053: begin
				if(in == 0) begin
					state<=7064;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=3175;
					out<=195;
				end
				if(in == 3) begin
					state<=5074;
					out<=196;
				end
				if(in == 4) begin
					state<=1176;
					out<=197;
				end
			end
			7054: begin
				if(in == 0) begin
					state<=7065;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=3176;
					out<=200;
				end
				if(in == 3) begin
					state<=5075;
					out<=201;
				end
				if(in == 4) begin
					state<=1177;
					out<=202;
				end
			end
			7055: begin
				if(in == 0) begin
					state<=7066;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=3177;
					out<=205;
				end
				if(in == 3) begin
					state<=5076;
					out<=206;
				end
				if(in == 4) begin
					state<=1178;
					out<=207;
				end
			end
			7056: begin
				if(in == 0) begin
					state<=7067;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=3178;
					out<=210;
				end
				if(in == 3) begin
					state<=5077;
					out<=211;
				end
				if(in == 4) begin
					state<=1179;
					out<=212;
				end
			end
			7057: begin
				if(in == 0) begin
					state<=7058;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=3169;
					out<=215;
				end
				if(in == 3) begin
					state<=5068;
					out<=216;
				end
				if(in == 4) begin
					state<=1170;
					out<=217;
				end
			end
			7058: begin
				if(in == 0) begin
					state<=7069;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=3180;
					out<=220;
				end
				if(in == 3) begin
					state<=5079;
					out<=221;
				end
				if(in == 4) begin
					state<=1181;
					out<=222;
				end
			end
			7059: begin
				if(in == 0) begin
					state<=7070;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=3181;
					out<=225;
				end
				if(in == 3) begin
					state<=5080;
					out<=226;
				end
				if(in == 4) begin
					state<=1182;
					out<=227;
				end
			end
			7060: begin
				if(in == 0) begin
					state<=7071;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=3182;
					out<=230;
				end
				if(in == 3) begin
					state<=5081;
					out<=231;
				end
				if(in == 4) begin
					state<=1183;
					out<=232;
				end
			end
			7061: begin
				if(in == 0) begin
					state<=7072;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=3183;
					out<=235;
				end
				if(in == 3) begin
					state<=5082;
					out<=236;
				end
				if(in == 4) begin
					state<=1184;
					out<=237;
				end
			end
			7062: begin
				if(in == 0) begin
					state<=7073;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=3184;
					out<=240;
				end
				if(in == 3) begin
					state<=5083;
					out<=241;
				end
				if(in == 4) begin
					state<=1185;
					out<=242;
				end
			end
			7063: begin
				if(in == 0) begin
					state<=7074;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=3185;
					out<=245;
				end
				if(in == 3) begin
					state<=5084;
					out<=246;
				end
				if(in == 4) begin
					state<=1186;
					out<=247;
				end
			end
			7064: begin
				if(in == 0) begin
					state<=7075;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=3186;
					out<=250;
				end
				if(in == 3) begin
					state<=5085;
					out<=251;
				end
				if(in == 4) begin
					state<=1187;
					out<=252;
				end
			end
			7065: begin
				if(in == 0) begin
					state<=7076;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=3187;
					out<=255;
				end
				if(in == 3) begin
					state<=5086;
					out<=0;
				end
				if(in == 4) begin
					state<=1188;
					out<=1;
				end
			end
			7066: begin
				if(in == 0) begin
					state<=7077;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=3188;
					out<=4;
				end
				if(in == 3) begin
					state<=5087;
					out<=5;
				end
				if(in == 4) begin
					state<=1189;
					out<=6;
				end
			end
			7067: begin
				if(in == 0) begin
					state<=7068;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=3179;
					out<=9;
				end
				if(in == 3) begin
					state<=5078;
					out<=10;
				end
				if(in == 4) begin
					state<=1180;
					out<=11;
				end
			end
			7068: begin
				if(in == 0) begin
					state<=7079;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=3190;
					out<=14;
				end
				if(in == 3) begin
					state<=5089;
					out<=15;
				end
				if(in == 4) begin
					state<=1191;
					out<=16;
				end
			end
			7069: begin
				if(in == 0) begin
					state<=7080;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=3191;
					out<=19;
				end
				if(in == 3) begin
					state<=5090;
					out<=20;
				end
				if(in == 4) begin
					state<=1192;
					out<=21;
				end
			end
			7070: begin
				if(in == 0) begin
					state<=7081;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=3192;
					out<=24;
				end
				if(in == 3) begin
					state<=5091;
					out<=25;
				end
				if(in == 4) begin
					state<=1193;
					out<=26;
				end
			end
			7071: begin
				if(in == 0) begin
					state<=7082;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=3193;
					out<=29;
				end
				if(in == 3) begin
					state<=5092;
					out<=30;
				end
				if(in == 4) begin
					state<=1194;
					out<=31;
				end
			end
			7072: begin
				if(in == 0) begin
					state<=7083;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=3194;
					out<=34;
				end
				if(in == 3) begin
					state<=5093;
					out<=35;
				end
				if(in == 4) begin
					state<=1195;
					out<=36;
				end
			end
			7073: begin
				if(in == 0) begin
					state<=7084;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=3195;
					out<=39;
				end
				if(in == 3) begin
					state<=5094;
					out<=40;
				end
				if(in == 4) begin
					state<=1196;
					out<=41;
				end
			end
			7074: begin
				if(in == 0) begin
					state<=7085;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=3196;
					out<=44;
				end
				if(in == 3) begin
					state<=5095;
					out<=45;
				end
				if(in == 4) begin
					state<=1197;
					out<=46;
				end
			end
			7075: begin
				if(in == 0) begin
					state<=7086;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=3197;
					out<=49;
				end
				if(in == 3) begin
					state<=5096;
					out<=50;
				end
				if(in == 4) begin
					state<=1198;
					out<=51;
				end
			end
			7076: begin
				if(in == 0) begin
					state<=7087;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=3198;
					out<=54;
				end
				if(in == 3) begin
					state<=5097;
					out<=55;
				end
				if(in == 4) begin
					state<=1199;
					out<=56;
				end
			end
			7077: begin
				if(in == 0) begin
					state<=7078;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=3189;
					out<=59;
				end
				if(in == 3) begin
					state<=5088;
					out<=60;
				end
				if(in == 4) begin
					state<=1190;
					out<=61;
				end
			end
			7078: begin
				if(in == 0) begin
					state<=7089;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=3200;
					out<=64;
				end
				if(in == 3) begin
					state<=5099;
					out<=65;
				end
				if(in == 4) begin
					state<=1201;
					out<=66;
				end
			end
			7079: begin
				if(in == 0) begin
					state<=7090;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=3201;
					out<=69;
				end
				if(in == 3) begin
					state<=5100;
					out<=70;
				end
				if(in == 4) begin
					state<=1202;
					out<=71;
				end
			end
			7080: begin
				if(in == 0) begin
					state<=7091;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=3202;
					out<=74;
				end
				if(in == 3) begin
					state<=5101;
					out<=75;
				end
				if(in == 4) begin
					state<=1203;
					out<=76;
				end
			end
			7081: begin
				if(in == 0) begin
					state<=7092;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=3203;
					out<=79;
				end
				if(in == 3) begin
					state<=5102;
					out<=80;
				end
				if(in == 4) begin
					state<=1204;
					out<=81;
				end
			end
			7082: begin
				if(in == 0) begin
					state<=7093;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=3204;
					out<=84;
				end
				if(in == 3) begin
					state<=5103;
					out<=85;
				end
				if(in == 4) begin
					state<=1205;
					out<=86;
				end
			end
			7083: begin
				if(in == 0) begin
					state<=7094;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=3205;
					out<=89;
				end
				if(in == 3) begin
					state<=5104;
					out<=90;
				end
				if(in == 4) begin
					state<=1206;
					out<=91;
				end
			end
			7084: begin
				if(in == 0) begin
					state<=7095;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=3206;
					out<=94;
				end
				if(in == 3) begin
					state<=5105;
					out<=95;
				end
				if(in == 4) begin
					state<=1207;
					out<=96;
				end
			end
			7085: begin
				if(in == 0) begin
					state<=7096;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=3207;
					out<=99;
				end
				if(in == 3) begin
					state<=5106;
					out<=100;
				end
				if(in == 4) begin
					state<=1208;
					out<=101;
				end
			end
			7086: begin
				if(in == 0) begin
					state<=7097;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=3208;
					out<=104;
				end
				if(in == 3) begin
					state<=5107;
					out<=105;
				end
				if(in == 4) begin
					state<=1209;
					out<=106;
				end
			end
			7087: begin
				if(in == 0) begin
					state<=7088;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=3199;
					out<=109;
				end
				if(in == 3) begin
					state<=5098;
					out<=110;
				end
				if(in == 4) begin
					state<=1200;
					out<=111;
				end
			end
			7088: begin
				if(in == 0) begin
					state<=7099;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=3210;
					out<=114;
				end
				if(in == 3) begin
					state<=5109;
					out<=115;
				end
				if(in == 4) begin
					state<=1211;
					out<=116;
				end
			end
			7089: begin
				if(in == 0) begin
					state<=7100;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=3211;
					out<=119;
				end
				if(in == 3) begin
					state<=5110;
					out<=120;
				end
				if(in == 4) begin
					state<=1212;
					out<=121;
				end
			end
			7090: begin
				if(in == 0) begin
					state<=7101;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=3212;
					out<=124;
				end
				if(in == 3) begin
					state<=5111;
					out<=125;
				end
				if(in == 4) begin
					state<=1213;
					out<=126;
				end
			end
			7091: begin
				if(in == 0) begin
					state<=7102;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=3213;
					out<=129;
				end
				if(in == 3) begin
					state<=5112;
					out<=130;
				end
				if(in == 4) begin
					state<=1214;
					out<=131;
				end
			end
			7092: begin
				if(in == 0) begin
					state<=7103;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=3214;
					out<=134;
				end
				if(in == 3) begin
					state<=5113;
					out<=135;
				end
				if(in == 4) begin
					state<=1215;
					out<=136;
				end
			end
			7093: begin
				if(in == 0) begin
					state<=7104;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=3215;
					out<=139;
				end
				if(in == 3) begin
					state<=5114;
					out<=140;
				end
				if(in == 4) begin
					state<=1216;
					out<=141;
				end
			end
			7094: begin
				if(in == 0) begin
					state<=7105;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=3216;
					out<=144;
				end
				if(in == 3) begin
					state<=5115;
					out<=145;
				end
				if(in == 4) begin
					state<=1217;
					out<=146;
				end
			end
			7095: begin
				if(in == 0) begin
					state<=7106;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=3217;
					out<=149;
				end
				if(in == 3) begin
					state<=5116;
					out<=150;
				end
				if(in == 4) begin
					state<=1218;
					out<=151;
				end
			end
			7096: begin
				if(in == 0) begin
					state<=7107;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=3218;
					out<=154;
				end
				if(in == 3) begin
					state<=5117;
					out<=155;
				end
				if(in == 4) begin
					state<=1219;
					out<=156;
				end
			end
			7097: begin
				if(in == 0) begin
					state<=7098;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=3209;
					out<=159;
				end
				if(in == 3) begin
					state<=5108;
					out<=160;
				end
				if(in == 4) begin
					state<=1210;
					out<=161;
				end
			end
			7098: begin
				if(in == 0) begin
					state<=7109;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=3220;
					out<=164;
				end
				if(in == 3) begin
					state<=5119;
					out<=165;
				end
				if(in == 4) begin
					state<=1221;
					out<=166;
				end
			end
			7099: begin
				if(in == 0) begin
					state<=7110;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=3221;
					out<=169;
				end
				if(in == 3) begin
					state<=5120;
					out<=170;
				end
				if(in == 4) begin
					state<=1222;
					out<=171;
				end
			end
			7100: begin
				if(in == 0) begin
					state<=7111;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=3222;
					out<=174;
				end
				if(in == 3) begin
					state<=5121;
					out<=175;
				end
				if(in == 4) begin
					state<=1223;
					out<=176;
				end
			end
			7101: begin
				if(in == 0) begin
					state<=7112;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=3223;
					out<=179;
				end
				if(in == 3) begin
					state<=5122;
					out<=180;
				end
				if(in == 4) begin
					state<=1224;
					out<=181;
				end
			end
			7102: begin
				if(in == 0) begin
					state<=7113;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=3224;
					out<=184;
				end
				if(in == 3) begin
					state<=5123;
					out<=185;
				end
				if(in == 4) begin
					state<=1225;
					out<=186;
				end
			end
			7103: begin
				if(in == 0) begin
					state<=7114;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=3225;
					out<=189;
				end
				if(in == 3) begin
					state<=5124;
					out<=190;
				end
				if(in == 4) begin
					state<=1226;
					out<=191;
				end
			end
			7104: begin
				if(in == 0) begin
					state<=7115;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=3226;
					out<=194;
				end
				if(in == 3) begin
					state<=5125;
					out<=195;
				end
				if(in == 4) begin
					state<=1227;
					out<=196;
				end
			end
			7105: begin
				if(in == 0) begin
					state<=7116;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=3227;
					out<=199;
				end
				if(in == 3) begin
					state<=5126;
					out<=200;
				end
				if(in == 4) begin
					state<=1228;
					out<=201;
				end
			end
			7106: begin
				if(in == 0) begin
					state<=7117;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=3228;
					out<=204;
				end
				if(in == 3) begin
					state<=5127;
					out<=205;
				end
				if(in == 4) begin
					state<=1229;
					out<=206;
				end
			end
			7107: begin
				if(in == 0) begin
					state<=7108;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=3219;
					out<=209;
				end
				if(in == 3) begin
					state<=5118;
					out<=210;
				end
				if(in == 4) begin
					state<=1220;
					out<=211;
				end
			end
			7108: begin
				if(in == 0) begin
					state<=6578;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=2689;
					out<=214;
				end
				if(in == 3) begin
					state<=4589;
					out<=215;
				end
				if(in == 4) begin
					state<=691;
					out<=216;
				end
			end
			7109: begin
				if(in == 0) begin
					state<=6579;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=2690;
					out<=219;
				end
				if(in == 3) begin
					state<=4590;
					out<=220;
				end
				if(in == 4) begin
					state<=692;
					out<=221;
				end
			end
			7110: begin
				if(in == 0) begin
					state<=6580;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=2691;
					out<=224;
				end
				if(in == 3) begin
					state<=4591;
					out<=225;
				end
				if(in == 4) begin
					state<=693;
					out<=226;
				end
			end
			7111: begin
				if(in == 0) begin
					state<=6581;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=2692;
					out<=229;
				end
				if(in == 3) begin
					state<=4592;
					out<=230;
				end
				if(in == 4) begin
					state<=694;
					out<=231;
				end
			end
			7112: begin
				if(in == 0) begin
					state<=6582;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=2693;
					out<=234;
				end
				if(in == 3) begin
					state<=4593;
					out<=235;
				end
				if(in == 4) begin
					state<=695;
					out<=236;
				end
			end
			7113: begin
				if(in == 0) begin
					state<=6583;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=2694;
					out<=239;
				end
				if(in == 3) begin
					state<=4594;
					out<=240;
				end
				if(in == 4) begin
					state<=696;
					out<=241;
				end
			end
			7114: begin
				if(in == 0) begin
					state<=6584;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=2695;
					out<=244;
				end
				if(in == 3) begin
					state<=4595;
					out<=245;
				end
				if(in == 4) begin
					state<=697;
					out<=246;
				end
			end
			7115: begin
				if(in == 0) begin
					state<=6585;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=2696;
					out<=249;
				end
				if(in == 3) begin
					state<=4596;
					out<=250;
				end
				if(in == 4) begin
					state<=698;
					out<=251;
				end
			end
			7116: begin
				if(in == 0) begin
					state<=6586;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=2697;
					out<=254;
				end
				if(in == 3) begin
					state<=4597;
					out<=255;
				end
				if(in == 4) begin
					state<=699;
					out<=0;
				end
			end
			7117: begin
				if(in == 0) begin
					state<=7118;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=3229;
					out<=3;
				end
				if(in == 3) begin
					state<=5128;
					out<=4;
				end
				if(in == 4) begin
					state<=1230;
					out<=5;
				end
			end
			7118: begin
				if(in == 0) begin
					state<=6588;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=2699;
					out<=8;
				end
				if(in == 3) begin
					state<=4599;
					out<=9;
				end
				if(in == 4) begin
					state<=701;
					out<=10;
				end
			end
			7119: begin
				if(in == 0) begin
					state<=7130;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=3241;
					out<=13;
				end
				if(in == 3) begin
					state<=5477;
					out<=14;
				end
				if(in == 4) begin
					state<=1588;
					out<=15;
				end
			end
			7120: begin
				if(in == 0) begin
					state<=7131;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=3242;
					out<=18;
				end
				if(in == 3) begin
					state<=5478;
					out<=19;
				end
				if(in == 4) begin
					state<=1589;
					out<=20;
				end
			end
			7121: begin
				if(in == 0) begin
					state<=7132;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=3243;
					out<=23;
				end
				if(in == 3) begin
					state<=5479;
					out<=24;
				end
				if(in == 4) begin
					state<=1590;
					out<=25;
				end
			end
			7122: begin
				if(in == 0) begin
					state<=7133;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=3244;
					out<=28;
				end
				if(in == 3) begin
					state<=5480;
					out<=29;
				end
				if(in == 4) begin
					state<=1591;
					out<=30;
				end
			end
			7123: begin
				if(in == 0) begin
					state<=7134;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=3245;
					out<=33;
				end
				if(in == 3) begin
					state<=5481;
					out<=34;
				end
				if(in == 4) begin
					state<=1592;
					out<=35;
				end
			end
			7124: begin
				if(in == 0) begin
					state<=7135;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=3246;
					out<=38;
				end
				if(in == 3) begin
					state<=5482;
					out<=39;
				end
				if(in == 4) begin
					state<=1593;
					out<=40;
				end
			end
			7125: begin
				if(in == 0) begin
					state<=7136;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=3247;
					out<=43;
				end
				if(in == 3) begin
					state<=5483;
					out<=44;
				end
				if(in == 4) begin
					state<=1594;
					out<=45;
				end
			end
			7126: begin
				if(in == 0) begin
					state<=7137;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=3248;
					out<=48;
				end
				if(in == 3) begin
					state<=5484;
					out<=49;
				end
				if(in == 4) begin
					state<=1595;
					out<=50;
				end
			end
			7127: begin
				if(in == 0) begin
					state<=7138;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=3249;
					out<=53;
				end
				if(in == 3) begin
					state<=5485;
					out<=54;
				end
				if(in == 4) begin
					state<=1596;
					out<=55;
				end
			end
			7128: begin
				if(in == 0) begin
					state<=7129;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=3240;
					out<=58;
				end
				if(in == 3) begin
					state<=5476;
					out<=59;
				end
				if(in == 4) begin
					state<=1587;
					out<=60;
				end
			end
			7129: begin
				if(in == 0) begin
					state<=7140;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=3251;
					out<=63;
				end
				if(in == 3) begin
					state<=5487;
					out<=64;
				end
				if(in == 4) begin
					state<=1598;
					out<=65;
				end
			end
			7130: begin
				if(in == 0) begin
					state<=7141;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=3252;
					out<=68;
				end
				if(in == 3) begin
					state<=5488;
					out<=69;
				end
				if(in == 4) begin
					state<=1599;
					out<=70;
				end
			end
			7131: begin
				if(in == 0) begin
					state<=7142;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=3253;
					out<=73;
				end
				if(in == 3) begin
					state<=5489;
					out<=74;
				end
				if(in == 4) begin
					state<=1600;
					out<=75;
				end
			end
			7132: begin
				if(in == 0) begin
					state<=7143;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=3254;
					out<=78;
				end
				if(in == 3) begin
					state<=5490;
					out<=79;
				end
				if(in == 4) begin
					state<=1601;
					out<=80;
				end
			end
			7133: begin
				if(in == 0) begin
					state<=7144;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=3255;
					out<=83;
				end
				if(in == 3) begin
					state<=5491;
					out<=84;
				end
				if(in == 4) begin
					state<=1602;
					out<=85;
				end
			end
			7134: begin
				if(in == 0) begin
					state<=7145;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=3256;
					out<=88;
				end
				if(in == 3) begin
					state<=5492;
					out<=89;
				end
				if(in == 4) begin
					state<=1603;
					out<=90;
				end
			end
			7135: begin
				if(in == 0) begin
					state<=7146;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=3257;
					out<=93;
				end
				if(in == 3) begin
					state<=5493;
					out<=94;
				end
				if(in == 4) begin
					state<=1604;
					out<=95;
				end
			end
			7136: begin
				if(in == 0) begin
					state<=7147;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=3258;
					out<=98;
				end
				if(in == 3) begin
					state<=5494;
					out<=99;
				end
				if(in == 4) begin
					state<=1605;
					out<=100;
				end
			end
			7137: begin
				if(in == 0) begin
					state<=7148;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=3259;
					out<=103;
				end
				if(in == 3) begin
					state<=5495;
					out<=104;
				end
				if(in == 4) begin
					state<=1606;
					out<=105;
				end
			end
			7138: begin
				if(in == 0) begin
					state<=7139;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=3250;
					out<=108;
				end
				if(in == 3) begin
					state<=5486;
					out<=109;
				end
				if(in == 4) begin
					state<=1597;
					out<=110;
				end
			end
			7139: begin
				if(in == 0) begin
					state<=6559;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=2670;
					out<=113;
				end
				if(in == 3) begin
					state<=4570;
					out<=114;
				end
				if(in == 4) begin
					state<=672;
					out<=115;
				end
			end
			7140: begin
				if(in == 0) begin
					state<=6560;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=2671;
					out<=118;
				end
				if(in == 3) begin
					state<=4571;
					out<=119;
				end
				if(in == 4) begin
					state<=673;
					out<=120;
				end
			end
			7141: begin
				if(in == 0) begin
					state<=6561;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=2672;
					out<=123;
				end
				if(in == 3) begin
					state<=4572;
					out<=124;
				end
				if(in == 4) begin
					state<=674;
					out<=125;
				end
			end
			7142: begin
				if(in == 0) begin
					state<=6562;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=2673;
					out<=128;
				end
				if(in == 3) begin
					state<=4573;
					out<=129;
				end
				if(in == 4) begin
					state<=675;
					out<=130;
				end
			end
			7143: begin
				if(in == 0) begin
					state<=6563;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=2674;
					out<=133;
				end
				if(in == 3) begin
					state<=4574;
					out<=134;
				end
				if(in == 4) begin
					state<=676;
					out<=135;
				end
			end
			7144: begin
				if(in == 0) begin
					state<=6564;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=2675;
					out<=138;
				end
				if(in == 3) begin
					state<=4575;
					out<=139;
				end
				if(in == 4) begin
					state<=677;
					out<=140;
				end
			end
			7145: begin
				if(in == 0) begin
					state<=6565;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=2676;
					out<=143;
				end
				if(in == 3) begin
					state<=4576;
					out<=144;
				end
				if(in == 4) begin
					state<=678;
					out<=145;
				end
			end
			7146: begin
				if(in == 0) begin
					state<=6566;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=2677;
					out<=148;
				end
				if(in == 3) begin
					state<=4577;
					out<=149;
				end
				if(in == 4) begin
					state<=679;
					out<=150;
				end
			end
			7147: begin
				if(in == 0) begin
					state<=6567;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=2678;
					out<=153;
				end
				if(in == 3) begin
					state<=4578;
					out<=154;
				end
				if(in == 4) begin
					state<=680;
					out<=155;
				end
			end
			7148: begin
				if(in == 0) begin
					state<=7149;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=3260;
					out<=158;
				end
				if(in == 3) begin
					state<=5496;
					out<=159;
				end
				if(in == 4) begin
					state<=1607;
					out<=160;
				end
			end
			7149: begin
				if(in == 0) begin
					state<=6569;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=2680;
					out<=163;
				end
				if(in == 3) begin
					state<=4580;
					out<=164;
				end
				if(in == 4) begin
					state<=682;
					out<=165;
				end
			end
			7150: begin
				if(in == 0) begin
					state<=7161;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=3272;
					out<=168;
				end
				if(in == 3) begin
					state<=5229;
					out<=169;
				end
				if(in == 4) begin
					state<=1340;
					out<=170;
				end
			end
			7151: begin
				if(in == 0) begin
					state<=7162;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=3273;
					out<=173;
				end
				if(in == 3) begin
					state<=5230;
					out<=174;
				end
				if(in == 4) begin
					state<=1341;
					out<=175;
				end
			end
			7152: begin
				if(in == 0) begin
					state<=7163;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=3274;
					out<=178;
				end
				if(in == 3) begin
					state<=5231;
					out<=179;
				end
				if(in == 4) begin
					state<=1342;
					out<=180;
				end
			end
			7153: begin
				if(in == 0) begin
					state<=7164;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=3275;
					out<=183;
				end
				if(in == 3) begin
					state<=5232;
					out<=184;
				end
				if(in == 4) begin
					state<=1343;
					out<=185;
				end
			end
			7154: begin
				if(in == 0) begin
					state<=7165;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=3276;
					out<=188;
				end
				if(in == 3) begin
					state<=5233;
					out<=189;
				end
				if(in == 4) begin
					state<=1344;
					out<=190;
				end
			end
			7155: begin
				if(in == 0) begin
					state<=7166;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=3277;
					out<=193;
				end
				if(in == 3) begin
					state<=5234;
					out<=194;
				end
				if(in == 4) begin
					state<=1345;
					out<=195;
				end
			end
			7156: begin
				if(in == 0) begin
					state<=7167;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=3278;
					out<=198;
				end
				if(in == 3) begin
					state<=5235;
					out<=199;
				end
				if(in == 4) begin
					state<=1346;
					out<=200;
				end
			end
			7157: begin
				if(in == 0) begin
					state<=7168;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=3279;
					out<=203;
				end
				if(in == 3) begin
					state<=5236;
					out<=204;
				end
				if(in == 4) begin
					state<=1347;
					out<=205;
				end
			end
			7158: begin
				if(in == 0) begin
					state<=7169;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=3280;
					out<=208;
				end
				if(in == 3) begin
					state<=5237;
					out<=209;
				end
				if(in == 4) begin
					state<=1348;
					out<=210;
				end
			end
			7159: begin
				if(in == 0) begin
					state<=7160;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=3271;
					out<=213;
				end
				if(in == 3) begin
					state<=5228;
					out<=214;
				end
				if(in == 4) begin
					state<=1339;
					out<=215;
				end
			end
			7160: begin
				if(in == 0) begin
					state<=7171;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=3282;
					out<=218;
				end
				if(in == 3) begin
					state<=5239;
					out<=219;
				end
				if(in == 4) begin
					state<=1350;
					out<=220;
				end
			end
			7161: begin
				if(in == 0) begin
					state<=7172;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=3283;
					out<=223;
				end
				if(in == 3) begin
					state<=5240;
					out<=224;
				end
				if(in == 4) begin
					state<=1351;
					out<=225;
				end
			end
			7162: begin
				if(in == 0) begin
					state<=7173;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=3284;
					out<=228;
				end
				if(in == 3) begin
					state<=5241;
					out<=229;
				end
				if(in == 4) begin
					state<=1352;
					out<=230;
				end
			end
			7163: begin
				if(in == 0) begin
					state<=7174;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=3285;
					out<=233;
				end
				if(in == 3) begin
					state<=5242;
					out<=234;
				end
				if(in == 4) begin
					state<=1353;
					out<=235;
				end
			end
			7164: begin
				if(in == 0) begin
					state<=7175;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=3286;
					out<=238;
				end
				if(in == 3) begin
					state<=5243;
					out<=239;
				end
				if(in == 4) begin
					state<=1354;
					out<=240;
				end
			end
			7165: begin
				if(in == 0) begin
					state<=7176;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=3287;
					out<=243;
				end
				if(in == 3) begin
					state<=5244;
					out<=244;
				end
				if(in == 4) begin
					state<=1355;
					out<=245;
				end
			end
			7166: begin
				if(in == 0) begin
					state<=7177;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=3288;
					out<=248;
				end
				if(in == 3) begin
					state<=5245;
					out<=249;
				end
				if(in == 4) begin
					state<=1356;
					out<=250;
				end
			end
			7167: begin
				if(in == 0) begin
					state<=7178;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=3289;
					out<=253;
				end
				if(in == 3) begin
					state<=5246;
					out<=254;
				end
				if(in == 4) begin
					state<=1357;
					out<=255;
				end
			end
			7168: begin
				if(in == 0) begin
					state<=7179;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=3290;
					out<=2;
				end
				if(in == 3) begin
					state<=5247;
					out<=3;
				end
				if(in == 4) begin
					state<=1358;
					out<=4;
				end
			end
			7169: begin
				if(in == 0) begin
					state<=7170;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=3281;
					out<=7;
				end
				if(in == 3) begin
					state<=5238;
					out<=8;
				end
				if(in == 4) begin
					state<=1349;
					out<=9;
				end
			end
			7170: begin
				if(in == 0) begin
					state<=5938;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=2049;
					out<=12;
				end
				if(in == 3) begin
					state<=3949;
					out<=13;
				end
				if(in == 4) begin
					state<=51;
					out<=14;
				end
			end
			7171: begin
				if(in == 0) begin
					state<=5939;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=2050;
					out<=17;
				end
				if(in == 3) begin
					state<=3950;
					out<=18;
				end
				if(in == 4) begin
					state<=52;
					out<=19;
				end
			end
			7172: begin
				if(in == 0) begin
					state<=5940;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=2051;
					out<=22;
				end
				if(in == 3) begin
					state<=3951;
					out<=23;
				end
				if(in == 4) begin
					state<=53;
					out<=24;
				end
			end
			7173: begin
				if(in == 0) begin
					state<=5941;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=2052;
					out<=27;
				end
				if(in == 3) begin
					state<=3952;
					out<=28;
				end
				if(in == 4) begin
					state<=54;
					out<=29;
				end
			end
			7174: begin
				if(in == 0) begin
					state<=5942;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=2053;
					out<=32;
				end
				if(in == 3) begin
					state<=3953;
					out<=33;
				end
				if(in == 4) begin
					state<=55;
					out<=34;
				end
			end
			7175: begin
				if(in == 0) begin
					state<=5943;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=2054;
					out<=37;
				end
				if(in == 3) begin
					state<=3954;
					out<=38;
				end
				if(in == 4) begin
					state<=56;
					out<=39;
				end
			end
			7176: begin
				if(in == 0) begin
					state<=5944;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=2055;
					out<=42;
				end
				if(in == 3) begin
					state<=3955;
					out<=43;
				end
				if(in == 4) begin
					state<=57;
					out<=44;
				end
			end
			7177: begin
				if(in == 0) begin
					state<=5945;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=2056;
					out<=47;
				end
				if(in == 3) begin
					state<=3956;
					out<=48;
				end
				if(in == 4) begin
					state<=58;
					out<=49;
				end
			end
			7178: begin
				if(in == 0) begin
					state<=5946;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=2057;
					out<=52;
				end
				if(in == 3) begin
					state<=3957;
					out<=53;
				end
				if(in == 4) begin
					state<=59;
					out<=54;
				end
			end
			7179: begin
				if(in == 0) begin
					state<=7180;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=3291;
					out<=57;
				end
				if(in == 3) begin
					state<=5248;
					out<=58;
				end
				if(in == 4) begin
					state<=1359;
					out<=59;
				end
			end
			7180: begin
				if(in == 0) begin
					state<=5948;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=2059;
					out<=62;
				end
				if(in == 3) begin
					state<=3959;
					out<=63;
				end
				if(in == 4) begin
					state<=61;
					out<=64;
				end
			end
			7181: begin
				if(in == 0) begin
					state<=7192;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=3303;
					out<=67;
				end
				if(in == 3) begin
					state<=5260;
					out<=68;
				end
				if(in == 4) begin
					state<=1371;
					out<=69;
				end
			end
			7182: begin
				if(in == 0) begin
					state<=7193;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=3304;
					out<=72;
				end
				if(in == 3) begin
					state<=5261;
					out<=73;
				end
				if(in == 4) begin
					state<=1372;
					out<=74;
				end
			end
			7183: begin
				if(in == 0) begin
					state<=7194;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=3305;
					out<=77;
				end
				if(in == 3) begin
					state<=5262;
					out<=78;
				end
				if(in == 4) begin
					state<=1373;
					out<=79;
				end
			end
			7184: begin
				if(in == 0) begin
					state<=7195;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=3306;
					out<=82;
				end
				if(in == 3) begin
					state<=5263;
					out<=83;
				end
				if(in == 4) begin
					state<=1374;
					out<=84;
				end
			end
			7185: begin
				if(in == 0) begin
					state<=7196;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=3307;
					out<=87;
				end
				if(in == 3) begin
					state<=5264;
					out<=88;
				end
				if(in == 4) begin
					state<=1375;
					out<=89;
				end
			end
			7186: begin
				if(in == 0) begin
					state<=7197;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=3308;
					out<=92;
				end
				if(in == 3) begin
					state<=5265;
					out<=93;
				end
				if(in == 4) begin
					state<=1376;
					out<=94;
				end
			end
			7187: begin
				if(in == 0) begin
					state<=7198;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=3309;
					out<=97;
				end
				if(in == 3) begin
					state<=5266;
					out<=98;
				end
				if(in == 4) begin
					state<=1377;
					out<=99;
				end
			end
			7188: begin
				if(in == 0) begin
					state<=7199;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=3310;
					out<=102;
				end
				if(in == 3) begin
					state<=5267;
					out<=103;
				end
				if(in == 4) begin
					state<=1378;
					out<=104;
				end
			end
			7189: begin
				if(in == 0) begin
					state<=7200;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=3311;
					out<=107;
				end
				if(in == 3) begin
					state<=5268;
					out<=108;
				end
				if(in == 4) begin
					state<=1379;
					out<=109;
				end
			end
			7190: begin
				if(in == 0) begin
					state<=7191;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=3302;
					out<=112;
				end
				if(in == 3) begin
					state<=5259;
					out<=113;
				end
				if(in == 4) begin
					state<=1370;
					out<=114;
				end
			end
			7191: begin
				if(in == 0) begin
					state<=7202;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=3313;
					out<=117;
				end
				if(in == 3) begin
					state<=5270;
					out<=118;
				end
				if(in == 4) begin
					state<=1381;
					out<=119;
				end
			end
			7192: begin
				if(in == 0) begin
					state<=7203;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=3314;
					out<=122;
				end
				if(in == 3) begin
					state<=5271;
					out<=123;
				end
				if(in == 4) begin
					state<=1382;
					out<=124;
				end
			end
			7193: begin
				if(in == 0) begin
					state<=7204;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=3315;
					out<=127;
				end
				if(in == 3) begin
					state<=5272;
					out<=128;
				end
				if(in == 4) begin
					state<=1383;
					out<=129;
				end
			end
			7194: begin
				if(in == 0) begin
					state<=7205;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=3316;
					out<=132;
				end
				if(in == 3) begin
					state<=5273;
					out<=133;
				end
				if(in == 4) begin
					state<=1384;
					out<=134;
				end
			end
			7195: begin
				if(in == 0) begin
					state<=7206;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=3317;
					out<=137;
				end
				if(in == 3) begin
					state<=5274;
					out<=138;
				end
				if(in == 4) begin
					state<=1385;
					out<=139;
				end
			end
			7196: begin
				if(in == 0) begin
					state<=7207;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=3318;
					out<=142;
				end
				if(in == 3) begin
					state<=5275;
					out<=143;
				end
				if(in == 4) begin
					state<=1386;
					out<=144;
				end
			end
			7197: begin
				if(in == 0) begin
					state<=7208;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=3319;
					out<=147;
				end
				if(in == 3) begin
					state<=5276;
					out<=148;
				end
				if(in == 4) begin
					state<=1387;
					out<=149;
				end
			end
			7198: begin
				if(in == 0) begin
					state<=7209;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=3320;
					out<=152;
				end
				if(in == 3) begin
					state<=5277;
					out<=153;
				end
				if(in == 4) begin
					state<=1388;
					out<=154;
				end
			end
			7199: begin
				if(in == 0) begin
					state<=7210;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=3321;
					out<=157;
				end
				if(in == 3) begin
					state<=5278;
					out<=158;
				end
				if(in == 4) begin
					state<=1389;
					out<=159;
				end
			end
			7200: begin
				if(in == 0) begin
					state<=7201;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=3312;
					out<=162;
				end
				if(in == 3) begin
					state<=5269;
					out<=163;
				end
				if(in == 4) begin
					state<=1380;
					out<=164;
				end
			end
			7201: begin
				if(in == 0) begin
					state<=6007;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=2118;
					out<=167;
				end
				if(in == 3) begin
					state<=4018;
					out<=168;
				end
				if(in == 4) begin
					state<=120;
					out<=169;
				end
			end
			7202: begin
				if(in == 0) begin
					state<=6008;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=2119;
					out<=172;
				end
				if(in == 3) begin
					state<=4019;
					out<=173;
				end
				if(in == 4) begin
					state<=121;
					out<=174;
				end
			end
			7203: begin
				if(in == 0) begin
					state<=6009;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=2120;
					out<=177;
				end
				if(in == 3) begin
					state<=4020;
					out<=178;
				end
				if(in == 4) begin
					state<=122;
					out<=179;
				end
			end
			7204: begin
				if(in == 0) begin
					state<=6010;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=2121;
					out<=182;
				end
				if(in == 3) begin
					state<=4021;
					out<=183;
				end
				if(in == 4) begin
					state<=123;
					out<=184;
				end
			end
			7205: begin
				if(in == 0) begin
					state<=6011;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=2122;
					out<=187;
				end
				if(in == 3) begin
					state<=4022;
					out<=188;
				end
				if(in == 4) begin
					state<=124;
					out<=189;
				end
			end
			7206: begin
				if(in == 0) begin
					state<=6012;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=2123;
					out<=192;
				end
				if(in == 3) begin
					state<=4023;
					out<=193;
				end
				if(in == 4) begin
					state<=125;
					out<=194;
				end
			end
			7207: begin
				if(in == 0) begin
					state<=6013;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=2124;
					out<=197;
				end
				if(in == 3) begin
					state<=4024;
					out<=198;
				end
				if(in == 4) begin
					state<=126;
					out<=199;
				end
			end
			7208: begin
				if(in == 0) begin
					state<=6014;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=2125;
					out<=202;
				end
				if(in == 3) begin
					state<=4025;
					out<=203;
				end
				if(in == 4) begin
					state<=127;
					out<=204;
				end
			end
			7209: begin
				if(in == 0) begin
					state<=6015;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=2126;
					out<=207;
				end
				if(in == 3) begin
					state<=4026;
					out<=208;
				end
				if(in == 4) begin
					state<=128;
					out<=209;
				end
			end
			7210: begin
				if(in == 0) begin
					state<=7211;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=3322;
					out<=212;
				end
				if(in == 3) begin
					state<=5279;
					out<=213;
				end
				if(in == 4) begin
					state<=1390;
					out<=214;
				end
			end
			7211: begin
				if(in == 0) begin
					state<=6017;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=2128;
					out<=217;
				end
				if(in == 3) begin
					state<=4028;
					out<=218;
				end
				if(in == 4) begin
					state<=130;
					out<=219;
				end
			end
			7212: begin
				if(in == 0) begin
					state<=7223;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=3334;
					out<=222;
				end
				if(in == 3) begin
					state<=5291;
					out<=223;
				end
				if(in == 4) begin
					state<=1402;
					out<=224;
				end
			end
			7213: begin
				if(in == 0) begin
					state<=7224;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=3335;
					out<=227;
				end
				if(in == 3) begin
					state<=5292;
					out<=228;
				end
				if(in == 4) begin
					state<=1403;
					out<=229;
				end
			end
			7214: begin
				if(in == 0) begin
					state<=7225;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=3336;
					out<=232;
				end
				if(in == 3) begin
					state<=5293;
					out<=233;
				end
				if(in == 4) begin
					state<=1404;
					out<=234;
				end
			end
			7215: begin
				if(in == 0) begin
					state<=7226;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=3337;
					out<=237;
				end
				if(in == 3) begin
					state<=5294;
					out<=238;
				end
				if(in == 4) begin
					state<=1405;
					out<=239;
				end
			end
			7216: begin
				if(in == 0) begin
					state<=7227;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=3338;
					out<=242;
				end
				if(in == 3) begin
					state<=5295;
					out<=243;
				end
				if(in == 4) begin
					state<=1406;
					out<=244;
				end
			end
			7217: begin
				if(in == 0) begin
					state<=7228;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=3339;
					out<=247;
				end
				if(in == 3) begin
					state<=5296;
					out<=248;
				end
				if(in == 4) begin
					state<=1407;
					out<=249;
				end
			end
			7218: begin
				if(in == 0) begin
					state<=7229;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=3340;
					out<=252;
				end
				if(in == 3) begin
					state<=5297;
					out<=253;
				end
				if(in == 4) begin
					state<=1408;
					out<=254;
				end
			end
			7219: begin
				if(in == 0) begin
					state<=7230;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=3341;
					out<=1;
				end
				if(in == 3) begin
					state<=5298;
					out<=2;
				end
				if(in == 4) begin
					state<=1409;
					out<=3;
				end
			end
			7220: begin
				if(in == 0) begin
					state<=7231;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=3342;
					out<=6;
				end
				if(in == 3) begin
					state<=5299;
					out<=7;
				end
				if(in == 4) begin
					state<=1410;
					out<=8;
				end
			end
			7221: begin
				if(in == 0) begin
					state<=7222;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=3333;
					out<=11;
				end
				if(in == 3) begin
					state<=5290;
					out<=12;
				end
				if(in == 4) begin
					state<=1401;
					out<=13;
				end
			end
			7222: begin
				if(in == 0) begin
					state<=7233;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=3344;
					out<=16;
				end
				if(in == 3) begin
					state<=5301;
					out<=17;
				end
				if(in == 4) begin
					state<=1412;
					out<=18;
				end
			end
			7223: begin
				if(in == 0) begin
					state<=7234;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=3345;
					out<=21;
				end
				if(in == 3) begin
					state<=5302;
					out<=22;
				end
				if(in == 4) begin
					state<=1413;
					out<=23;
				end
			end
			7224: begin
				if(in == 0) begin
					state<=7235;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=3346;
					out<=26;
				end
				if(in == 3) begin
					state<=5303;
					out<=27;
				end
				if(in == 4) begin
					state<=1414;
					out<=28;
				end
			end
			7225: begin
				if(in == 0) begin
					state<=7236;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=3347;
					out<=31;
				end
				if(in == 3) begin
					state<=5304;
					out<=32;
				end
				if(in == 4) begin
					state<=1415;
					out<=33;
				end
			end
			7226: begin
				if(in == 0) begin
					state<=7237;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=3348;
					out<=36;
				end
				if(in == 3) begin
					state<=5305;
					out<=37;
				end
				if(in == 4) begin
					state<=1416;
					out<=38;
				end
			end
			7227: begin
				if(in == 0) begin
					state<=7238;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=3349;
					out<=41;
				end
				if(in == 3) begin
					state<=5306;
					out<=42;
				end
				if(in == 4) begin
					state<=1417;
					out<=43;
				end
			end
			7228: begin
				if(in == 0) begin
					state<=7239;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=3350;
					out<=46;
				end
				if(in == 3) begin
					state<=5307;
					out<=47;
				end
				if(in == 4) begin
					state<=1418;
					out<=48;
				end
			end
			7229: begin
				if(in == 0) begin
					state<=7240;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=3351;
					out<=51;
				end
				if(in == 3) begin
					state<=5308;
					out<=52;
				end
				if(in == 4) begin
					state<=1419;
					out<=53;
				end
			end
			7230: begin
				if(in == 0) begin
					state<=7241;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=3352;
					out<=56;
				end
				if(in == 3) begin
					state<=5309;
					out<=57;
				end
				if(in == 4) begin
					state<=1420;
					out<=58;
				end
			end
			7231: begin
				if(in == 0) begin
					state<=7232;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=3343;
					out<=61;
				end
				if(in == 3) begin
					state<=5300;
					out<=62;
				end
				if(in == 4) begin
					state<=1411;
					out<=63;
				end
			end
			7232: begin
				if(in == 0) begin
					state<=6076;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=2187;
					out<=66;
				end
				if(in == 3) begin
					state<=4087;
					out<=67;
				end
				if(in == 4) begin
					state<=189;
					out<=68;
				end
			end
			7233: begin
				if(in == 0) begin
					state<=6077;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=2188;
					out<=71;
				end
				if(in == 3) begin
					state<=4088;
					out<=72;
				end
				if(in == 4) begin
					state<=190;
					out<=73;
				end
			end
			7234: begin
				if(in == 0) begin
					state<=6078;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=2189;
					out<=76;
				end
				if(in == 3) begin
					state<=4089;
					out<=77;
				end
				if(in == 4) begin
					state<=191;
					out<=78;
				end
			end
			7235: begin
				if(in == 0) begin
					state<=6079;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=2190;
					out<=81;
				end
				if(in == 3) begin
					state<=4090;
					out<=82;
				end
				if(in == 4) begin
					state<=192;
					out<=83;
				end
			end
			7236: begin
				if(in == 0) begin
					state<=6080;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=2191;
					out<=86;
				end
				if(in == 3) begin
					state<=4091;
					out<=87;
				end
				if(in == 4) begin
					state<=193;
					out<=88;
				end
			end
			7237: begin
				if(in == 0) begin
					state<=6081;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=2192;
					out<=91;
				end
				if(in == 3) begin
					state<=4092;
					out<=92;
				end
				if(in == 4) begin
					state<=194;
					out<=93;
				end
			end
			7238: begin
				if(in == 0) begin
					state<=6082;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=2193;
					out<=96;
				end
				if(in == 3) begin
					state<=4093;
					out<=97;
				end
				if(in == 4) begin
					state<=195;
					out<=98;
				end
			end
			7239: begin
				if(in == 0) begin
					state<=6083;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=2194;
					out<=101;
				end
				if(in == 3) begin
					state<=4094;
					out<=102;
				end
				if(in == 4) begin
					state<=196;
					out<=103;
				end
			end
			7240: begin
				if(in == 0) begin
					state<=6084;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=2195;
					out<=106;
				end
				if(in == 3) begin
					state<=4095;
					out<=107;
				end
				if(in == 4) begin
					state<=197;
					out<=108;
				end
			end
			7241: begin
				if(in == 0) begin
					state<=7242;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=3353;
					out<=111;
				end
				if(in == 3) begin
					state<=5310;
					out<=112;
				end
				if(in == 4) begin
					state<=1421;
					out<=113;
				end
			end
			7242: begin
				if(in == 0) begin
					state<=6086;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=2197;
					out<=116;
				end
				if(in == 3) begin
					state<=4097;
					out<=117;
				end
				if(in == 4) begin
					state<=199;
					out<=118;
				end
			end
			7243: begin
				if(in == 0) begin
					state<=7254;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=3365;
					out<=121;
				end
				if(in == 3) begin
					state<=5322;
					out<=122;
				end
				if(in == 4) begin
					state<=1433;
					out<=123;
				end
			end
			7244: begin
				if(in == 0) begin
					state<=7255;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=3366;
					out<=126;
				end
				if(in == 3) begin
					state<=5323;
					out<=127;
				end
				if(in == 4) begin
					state<=1434;
					out<=128;
				end
			end
			7245: begin
				if(in == 0) begin
					state<=7256;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=3367;
					out<=131;
				end
				if(in == 3) begin
					state<=5324;
					out<=132;
				end
				if(in == 4) begin
					state<=1435;
					out<=133;
				end
			end
			7246: begin
				if(in == 0) begin
					state<=7257;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=3368;
					out<=136;
				end
				if(in == 3) begin
					state<=5325;
					out<=137;
				end
				if(in == 4) begin
					state<=1436;
					out<=138;
				end
			end
			7247: begin
				if(in == 0) begin
					state<=7258;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=3369;
					out<=141;
				end
				if(in == 3) begin
					state<=5326;
					out<=142;
				end
				if(in == 4) begin
					state<=1437;
					out<=143;
				end
			end
			7248: begin
				if(in == 0) begin
					state<=7259;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=3370;
					out<=146;
				end
				if(in == 3) begin
					state<=5327;
					out<=147;
				end
				if(in == 4) begin
					state<=1438;
					out<=148;
				end
			end
			7249: begin
				if(in == 0) begin
					state<=7260;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=3371;
					out<=151;
				end
				if(in == 3) begin
					state<=5328;
					out<=152;
				end
				if(in == 4) begin
					state<=1439;
					out<=153;
				end
			end
			7250: begin
				if(in == 0) begin
					state<=7261;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=3372;
					out<=156;
				end
				if(in == 3) begin
					state<=5329;
					out<=157;
				end
				if(in == 4) begin
					state<=1440;
					out<=158;
				end
			end
			7251: begin
				if(in == 0) begin
					state<=7262;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=3373;
					out<=161;
				end
				if(in == 3) begin
					state<=5330;
					out<=162;
				end
				if(in == 4) begin
					state<=1441;
					out<=163;
				end
			end
			7252: begin
				if(in == 0) begin
					state<=7253;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=3364;
					out<=166;
				end
				if(in == 3) begin
					state<=5321;
					out<=167;
				end
				if(in == 4) begin
					state<=1432;
					out<=168;
				end
			end
			7253: begin
				if(in == 0) begin
					state<=7264;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=3375;
					out<=171;
				end
				if(in == 3) begin
					state<=5332;
					out<=172;
				end
				if(in == 4) begin
					state<=1443;
					out<=173;
				end
			end
			7254: begin
				if(in == 0) begin
					state<=7265;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=3376;
					out<=176;
				end
				if(in == 3) begin
					state<=5333;
					out<=177;
				end
				if(in == 4) begin
					state<=1444;
					out<=178;
				end
			end
			7255: begin
				if(in == 0) begin
					state<=7266;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=3377;
					out<=181;
				end
				if(in == 3) begin
					state<=5334;
					out<=182;
				end
				if(in == 4) begin
					state<=1445;
					out<=183;
				end
			end
			7256: begin
				if(in == 0) begin
					state<=7267;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=3378;
					out<=186;
				end
				if(in == 3) begin
					state<=5335;
					out<=187;
				end
				if(in == 4) begin
					state<=1446;
					out<=188;
				end
			end
			7257: begin
				if(in == 0) begin
					state<=7268;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=3379;
					out<=191;
				end
				if(in == 3) begin
					state<=5336;
					out<=192;
				end
				if(in == 4) begin
					state<=1447;
					out<=193;
				end
			end
			7258: begin
				if(in == 0) begin
					state<=7269;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=3380;
					out<=196;
				end
				if(in == 3) begin
					state<=5337;
					out<=197;
				end
				if(in == 4) begin
					state<=1448;
					out<=198;
				end
			end
			7259: begin
				if(in == 0) begin
					state<=7270;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=3381;
					out<=201;
				end
				if(in == 3) begin
					state<=5338;
					out<=202;
				end
				if(in == 4) begin
					state<=1449;
					out<=203;
				end
			end
			7260: begin
				if(in == 0) begin
					state<=7271;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=3382;
					out<=206;
				end
				if(in == 3) begin
					state<=5339;
					out<=207;
				end
				if(in == 4) begin
					state<=1450;
					out<=208;
				end
			end
			7261: begin
				if(in == 0) begin
					state<=7272;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=3383;
					out<=211;
				end
				if(in == 3) begin
					state<=5340;
					out<=212;
				end
				if(in == 4) begin
					state<=1451;
					out<=213;
				end
			end
			7262: begin
				if(in == 0) begin
					state<=7263;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=3374;
					out<=216;
				end
				if(in == 3) begin
					state<=5331;
					out<=217;
				end
				if(in == 4) begin
					state<=1442;
					out<=218;
				end
			end
			7263: begin
				if(in == 0) begin
					state<=6145;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=2256;
					out<=221;
				end
				if(in == 3) begin
					state<=4156;
					out<=222;
				end
				if(in == 4) begin
					state<=258;
					out<=223;
				end
			end
			7264: begin
				if(in == 0) begin
					state<=6146;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=2257;
					out<=226;
				end
				if(in == 3) begin
					state<=4157;
					out<=227;
				end
				if(in == 4) begin
					state<=259;
					out<=228;
				end
			end
			7265: begin
				if(in == 0) begin
					state<=6147;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=2258;
					out<=231;
				end
				if(in == 3) begin
					state<=4158;
					out<=232;
				end
				if(in == 4) begin
					state<=260;
					out<=233;
				end
			end
			7266: begin
				if(in == 0) begin
					state<=6148;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=2259;
					out<=236;
				end
				if(in == 3) begin
					state<=4159;
					out<=237;
				end
				if(in == 4) begin
					state<=261;
					out<=238;
				end
			end
			7267: begin
				if(in == 0) begin
					state<=6149;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=2260;
					out<=241;
				end
				if(in == 3) begin
					state<=4160;
					out<=242;
				end
				if(in == 4) begin
					state<=262;
					out<=243;
				end
			end
			7268: begin
				if(in == 0) begin
					state<=6150;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=2261;
					out<=246;
				end
				if(in == 3) begin
					state<=4161;
					out<=247;
				end
				if(in == 4) begin
					state<=263;
					out<=248;
				end
			end
			7269: begin
				if(in == 0) begin
					state<=6151;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=2262;
					out<=251;
				end
				if(in == 3) begin
					state<=4162;
					out<=252;
				end
				if(in == 4) begin
					state<=264;
					out<=253;
				end
			end
			7270: begin
				if(in == 0) begin
					state<=6152;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=2263;
					out<=0;
				end
				if(in == 3) begin
					state<=4163;
					out<=1;
				end
				if(in == 4) begin
					state<=265;
					out<=2;
				end
			end
			7271: begin
				if(in == 0) begin
					state<=6153;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=2264;
					out<=5;
				end
				if(in == 3) begin
					state<=4164;
					out<=6;
				end
				if(in == 4) begin
					state<=266;
					out<=7;
				end
			end
			7272: begin
				if(in == 0) begin
					state<=7273;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=3384;
					out<=10;
				end
				if(in == 3) begin
					state<=5341;
					out<=11;
				end
				if(in == 4) begin
					state<=1452;
					out<=12;
				end
			end
			7273: begin
				if(in == 0) begin
					state<=6155;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=2266;
					out<=15;
				end
				if(in == 3) begin
					state<=4166;
					out<=16;
				end
				if(in == 4) begin
					state<=268;
					out<=17;
				end
			end
			7274: begin
				if(in == 0) begin
					state<=7285;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=3396;
					out<=20;
				end
				if(in == 3) begin
					state<=4908;
					out<=21;
				end
				if(in == 4) begin
					state<=1010;
					out<=22;
				end
			end
			7275: begin
				if(in == 0) begin
					state<=7286;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=3397;
					out<=25;
				end
				if(in == 3) begin
					state<=4909;
					out<=26;
				end
				if(in == 4) begin
					state<=1011;
					out<=27;
				end
			end
			7276: begin
				if(in == 0) begin
					state<=7287;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=3398;
					out<=30;
				end
				if(in == 3) begin
					state<=4910;
					out<=31;
				end
				if(in == 4) begin
					state<=1012;
					out<=32;
				end
			end
			7277: begin
				if(in == 0) begin
					state<=7288;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=3399;
					out<=35;
				end
				if(in == 3) begin
					state<=4911;
					out<=36;
				end
				if(in == 4) begin
					state<=1013;
					out<=37;
				end
			end
			7278: begin
				if(in == 0) begin
					state<=7289;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=3400;
					out<=40;
				end
				if(in == 3) begin
					state<=4912;
					out<=41;
				end
				if(in == 4) begin
					state<=1014;
					out<=42;
				end
			end
			7279: begin
				if(in == 0) begin
					state<=7290;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=3401;
					out<=45;
				end
				if(in == 3) begin
					state<=4913;
					out<=46;
				end
				if(in == 4) begin
					state<=1015;
					out<=47;
				end
			end
			7280: begin
				if(in == 0) begin
					state<=7291;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=3402;
					out<=50;
				end
				if(in == 3) begin
					state<=4914;
					out<=51;
				end
				if(in == 4) begin
					state<=1016;
					out<=52;
				end
			end
			7281: begin
				if(in == 0) begin
					state<=7292;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=3403;
					out<=55;
				end
				if(in == 3) begin
					state<=4915;
					out<=56;
				end
				if(in == 4) begin
					state<=1017;
					out<=57;
				end
			end
			7282: begin
				if(in == 0) begin
					state<=7293;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=3404;
					out<=60;
				end
				if(in == 3) begin
					state<=4916;
					out<=61;
				end
				if(in == 4) begin
					state<=1018;
					out<=62;
				end
			end
			7283: begin
				if(in == 0) begin
					state<=7284;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=3395;
					out<=65;
				end
				if(in == 3) begin
					state<=4907;
					out<=66;
				end
				if(in == 4) begin
					state<=1009;
					out<=67;
				end
			end
			7284: begin
				if(in == 0) begin
					state<=7295;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=3406;
					out<=70;
				end
				if(in == 3) begin
					state<=4918;
					out<=71;
				end
				if(in == 4) begin
					state<=1020;
					out<=72;
				end
			end
			7285: begin
				if(in == 0) begin
					state<=7296;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=3407;
					out<=75;
				end
				if(in == 3) begin
					state<=4919;
					out<=76;
				end
				if(in == 4) begin
					state<=1021;
					out<=77;
				end
			end
			7286: begin
				if(in == 0) begin
					state<=7297;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=3408;
					out<=80;
				end
				if(in == 3) begin
					state<=4920;
					out<=81;
				end
				if(in == 4) begin
					state<=1022;
					out<=82;
				end
			end
			7287: begin
				if(in == 0) begin
					state<=7298;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=3409;
					out<=85;
				end
				if(in == 3) begin
					state<=4921;
					out<=86;
				end
				if(in == 4) begin
					state<=1023;
					out<=87;
				end
			end
			7288: begin
				if(in == 0) begin
					state<=7299;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=3410;
					out<=90;
				end
				if(in == 3) begin
					state<=4922;
					out<=91;
				end
				if(in == 4) begin
					state<=1024;
					out<=92;
				end
			end
			7289: begin
				if(in == 0) begin
					state<=7300;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=3411;
					out<=95;
				end
				if(in == 3) begin
					state<=4923;
					out<=96;
				end
				if(in == 4) begin
					state<=1025;
					out<=97;
				end
			end
			7290: begin
				if(in == 0) begin
					state<=7301;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=3412;
					out<=100;
				end
				if(in == 3) begin
					state<=4924;
					out<=101;
				end
				if(in == 4) begin
					state<=1026;
					out<=102;
				end
			end
			7291: begin
				if(in == 0) begin
					state<=7302;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=3413;
					out<=105;
				end
				if(in == 3) begin
					state<=4925;
					out<=106;
				end
				if(in == 4) begin
					state<=1027;
					out<=107;
				end
			end
			7292: begin
				if(in == 0) begin
					state<=7303;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=3414;
					out<=110;
				end
				if(in == 3) begin
					state<=4926;
					out<=111;
				end
				if(in == 4) begin
					state<=1028;
					out<=112;
				end
			end
			7293: begin
				if(in == 0) begin
					state<=7294;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=3405;
					out<=115;
				end
				if(in == 3) begin
					state<=4917;
					out<=116;
				end
				if(in == 4) begin
					state<=1019;
					out<=117;
				end
			end
			7294: begin
				if(in == 0) begin
					state<=6283;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=2394;
					out<=120;
				end
				if(in == 3) begin
					state<=4294;
					out<=121;
				end
				if(in == 4) begin
					state<=396;
					out<=122;
				end
			end
			7295: begin
				if(in == 0) begin
					state<=6284;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=2395;
					out<=125;
				end
				if(in == 3) begin
					state<=4295;
					out<=126;
				end
				if(in == 4) begin
					state<=397;
					out<=127;
				end
			end
			7296: begin
				if(in == 0) begin
					state<=6285;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=2396;
					out<=130;
				end
				if(in == 3) begin
					state<=4296;
					out<=131;
				end
				if(in == 4) begin
					state<=398;
					out<=132;
				end
			end
			7297: begin
				if(in == 0) begin
					state<=6286;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=2397;
					out<=135;
				end
				if(in == 3) begin
					state<=4297;
					out<=136;
				end
				if(in == 4) begin
					state<=399;
					out<=137;
				end
			end
			7298: begin
				if(in == 0) begin
					state<=6287;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=2398;
					out<=140;
				end
				if(in == 3) begin
					state<=4298;
					out<=141;
				end
				if(in == 4) begin
					state<=400;
					out<=142;
				end
			end
			7299: begin
				if(in == 0) begin
					state<=6288;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=2399;
					out<=145;
				end
				if(in == 3) begin
					state<=4299;
					out<=146;
				end
				if(in == 4) begin
					state<=401;
					out<=147;
				end
			end
			7300: begin
				if(in == 0) begin
					state<=6289;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=2400;
					out<=150;
				end
				if(in == 3) begin
					state<=4300;
					out<=151;
				end
				if(in == 4) begin
					state<=402;
					out<=152;
				end
			end
			7301: begin
				if(in == 0) begin
					state<=6290;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=2401;
					out<=155;
				end
				if(in == 3) begin
					state<=4301;
					out<=156;
				end
				if(in == 4) begin
					state<=403;
					out<=157;
				end
			end
			7302: begin
				if(in == 0) begin
					state<=6291;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=2402;
					out<=160;
				end
				if(in == 3) begin
					state<=4302;
					out<=161;
				end
				if(in == 4) begin
					state<=404;
					out<=162;
				end
			end
			7303: begin
				if(in == 0) begin
					state<=7304;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=3415;
					out<=165;
				end
				if(in == 3) begin
					state<=4927;
					out<=166;
				end
				if(in == 4) begin
					state<=1029;
					out<=167;
				end
			end
			7304: begin
				if(in == 0) begin
					state<=6293;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=2404;
					out<=170;
				end
				if(in == 3) begin
					state<=4304;
					out<=171;
				end
				if(in == 4) begin
					state<=406;
					out<=172;
				end
			end
			7305: begin
				if(in == 0) begin
					state<=7316;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=3427;
					out<=175;
				end
				if(in == 3) begin
					state<=5384;
					out<=176;
				end
				if(in == 4) begin
					state<=1495;
					out<=177;
				end
			end
			7306: begin
				if(in == 0) begin
					state<=7317;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=3428;
					out<=180;
				end
				if(in == 3) begin
					state<=5385;
					out<=181;
				end
				if(in == 4) begin
					state<=1496;
					out<=182;
				end
			end
			7307: begin
				if(in == 0) begin
					state<=7318;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=3429;
					out<=185;
				end
				if(in == 3) begin
					state<=5386;
					out<=186;
				end
				if(in == 4) begin
					state<=1497;
					out<=187;
				end
			end
			7308: begin
				if(in == 0) begin
					state<=7319;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=3430;
					out<=190;
				end
				if(in == 3) begin
					state<=5387;
					out<=191;
				end
				if(in == 4) begin
					state<=1498;
					out<=192;
				end
			end
			7309: begin
				if(in == 0) begin
					state<=7320;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=3431;
					out<=195;
				end
				if(in == 3) begin
					state<=5388;
					out<=196;
				end
				if(in == 4) begin
					state<=1499;
					out<=197;
				end
			end
			7310: begin
				if(in == 0) begin
					state<=7321;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=3432;
					out<=200;
				end
				if(in == 3) begin
					state<=5389;
					out<=201;
				end
				if(in == 4) begin
					state<=1500;
					out<=202;
				end
			end
			7311: begin
				if(in == 0) begin
					state<=7322;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=3433;
					out<=205;
				end
				if(in == 3) begin
					state<=5390;
					out<=206;
				end
				if(in == 4) begin
					state<=1501;
					out<=207;
				end
			end
			7312: begin
				if(in == 0) begin
					state<=7323;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=3434;
					out<=210;
				end
				if(in == 3) begin
					state<=5391;
					out<=211;
				end
				if(in == 4) begin
					state<=1502;
					out<=212;
				end
			end
			7313: begin
				if(in == 0) begin
					state<=7324;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=3435;
					out<=215;
				end
				if(in == 3) begin
					state<=5392;
					out<=216;
				end
				if(in == 4) begin
					state<=1503;
					out<=217;
				end
			end
			7314: begin
				if(in == 0) begin
					state<=7315;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=3426;
					out<=220;
				end
				if(in == 3) begin
					state<=5383;
					out<=221;
				end
				if(in == 4) begin
					state<=1494;
					out<=222;
				end
			end
			7315: begin
				if(in == 0) begin
					state<=7326;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=3437;
					out<=225;
				end
				if(in == 3) begin
					state<=5394;
					out<=226;
				end
				if(in == 4) begin
					state<=1505;
					out<=227;
				end
			end
			7316: begin
				if(in == 0) begin
					state<=7327;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=3438;
					out<=230;
				end
				if(in == 3) begin
					state<=5395;
					out<=231;
				end
				if(in == 4) begin
					state<=1506;
					out<=232;
				end
			end
			7317: begin
				if(in == 0) begin
					state<=7328;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=3439;
					out<=235;
				end
				if(in == 3) begin
					state<=5396;
					out<=236;
				end
				if(in == 4) begin
					state<=1507;
					out<=237;
				end
			end
			7318: begin
				if(in == 0) begin
					state<=7329;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=3440;
					out<=240;
				end
				if(in == 3) begin
					state<=5397;
					out<=241;
				end
				if(in == 4) begin
					state<=1508;
					out<=242;
				end
			end
			7319: begin
				if(in == 0) begin
					state<=7330;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=3441;
					out<=245;
				end
				if(in == 3) begin
					state<=5398;
					out<=246;
				end
				if(in == 4) begin
					state<=1509;
					out<=247;
				end
			end
			7320: begin
				if(in == 0) begin
					state<=7331;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=3442;
					out<=250;
				end
				if(in == 3) begin
					state<=5399;
					out<=251;
				end
				if(in == 4) begin
					state<=1510;
					out<=252;
				end
			end
			7321: begin
				if(in == 0) begin
					state<=7332;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=3443;
					out<=255;
				end
				if(in == 3) begin
					state<=5400;
					out<=0;
				end
				if(in == 4) begin
					state<=1511;
					out<=1;
				end
			end
			7322: begin
				if(in == 0) begin
					state<=7333;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=3444;
					out<=4;
				end
				if(in == 3) begin
					state<=5401;
					out<=5;
				end
				if(in == 4) begin
					state<=1512;
					out<=6;
				end
			end
			7323: begin
				if(in == 0) begin
					state<=7334;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=3445;
					out<=9;
				end
				if(in == 3) begin
					state<=5402;
					out<=10;
				end
				if(in == 4) begin
					state<=1513;
					out<=11;
				end
			end
			7324: begin
				if(in == 0) begin
					state<=7325;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=3436;
					out<=14;
				end
				if(in == 3) begin
					state<=5393;
					out<=15;
				end
				if(in == 4) begin
					state<=1504;
					out<=16;
				end
			end
			7325: begin
				if(in == 0) begin
					state<=6352;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=2463;
					out<=19;
				end
				if(in == 3) begin
					state<=4363;
					out<=20;
				end
				if(in == 4) begin
					state<=465;
					out<=21;
				end
			end
			7326: begin
				if(in == 0) begin
					state<=6353;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=2464;
					out<=24;
				end
				if(in == 3) begin
					state<=4364;
					out<=25;
				end
				if(in == 4) begin
					state<=466;
					out<=26;
				end
			end
			7327: begin
				if(in == 0) begin
					state<=6354;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=2465;
					out<=29;
				end
				if(in == 3) begin
					state<=4365;
					out<=30;
				end
				if(in == 4) begin
					state<=467;
					out<=31;
				end
			end
			7328: begin
				if(in == 0) begin
					state<=6355;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=2466;
					out<=34;
				end
				if(in == 3) begin
					state<=4366;
					out<=35;
				end
				if(in == 4) begin
					state<=468;
					out<=36;
				end
			end
			7329: begin
				if(in == 0) begin
					state<=6356;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=2467;
					out<=39;
				end
				if(in == 3) begin
					state<=4367;
					out<=40;
				end
				if(in == 4) begin
					state<=469;
					out<=41;
				end
			end
			7330: begin
				if(in == 0) begin
					state<=6357;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=2468;
					out<=44;
				end
				if(in == 3) begin
					state<=4368;
					out<=45;
				end
				if(in == 4) begin
					state<=470;
					out<=46;
				end
			end
			7331: begin
				if(in == 0) begin
					state<=6358;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=2469;
					out<=49;
				end
				if(in == 3) begin
					state<=4369;
					out<=50;
				end
				if(in == 4) begin
					state<=471;
					out<=51;
				end
			end
			7332: begin
				if(in == 0) begin
					state<=6359;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=2470;
					out<=54;
				end
				if(in == 3) begin
					state<=4370;
					out<=55;
				end
				if(in == 4) begin
					state<=472;
					out<=56;
				end
			end
			7333: begin
				if(in == 0) begin
					state<=6360;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=2471;
					out<=59;
				end
				if(in == 3) begin
					state<=4371;
					out<=60;
				end
				if(in == 4) begin
					state<=473;
					out<=61;
				end
			end
			7334: begin
				if(in == 0) begin
					state<=7335;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=3446;
					out<=64;
				end
				if(in == 3) begin
					state<=5403;
					out<=65;
				end
				if(in == 4) begin
					state<=1514;
					out<=66;
				end
			end
			7335: begin
				if(in == 0) begin
					state<=6362;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=2473;
					out<=69;
				end
				if(in == 3) begin
					state<=4373;
					out<=70;
				end
				if(in == 4) begin
					state<=475;
					out<=71;
				end
			end
			7336: begin
				if(in == 0) begin
					state<=7347;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=3458;
					out<=74;
				end
				if(in == 3) begin
					state<=5415;
					out<=75;
				end
				if(in == 4) begin
					state<=1526;
					out<=76;
				end
			end
			7337: begin
				if(in == 0) begin
					state<=7348;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=3459;
					out<=79;
				end
				if(in == 3) begin
					state<=5416;
					out<=80;
				end
				if(in == 4) begin
					state<=1527;
					out<=81;
				end
			end
			7338: begin
				if(in == 0) begin
					state<=7349;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=3460;
					out<=84;
				end
				if(in == 3) begin
					state<=5417;
					out<=85;
				end
				if(in == 4) begin
					state<=1528;
					out<=86;
				end
			end
			7339: begin
				if(in == 0) begin
					state<=7350;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=3461;
					out<=89;
				end
				if(in == 3) begin
					state<=5418;
					out<=90;
				end
				if(in == 4) begin
					state<=1529;
					out<=91;
				end
			end
			7340: begin
				if(in == 0) begin
					state<=7351;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=3462;
					out<=94;
				end
				if(in == 3) begin
					state<=5419;
					out<=95;
				end
				if(in == 4) begin
					state<=1530;
					out<=96;
				end
			end
			7341: begin
				if(in == 0) begin
					state<=7352;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=3463;
					out<=99;
				end
				if(in == 3) begin
					state<=5420;
					out<=100;
				end
				if(in == 4) begin
					state<=1531;
					out<=101;
				end
			end
			7342: begin
				if(in == 0) begin
					state<=7353;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=3464;
					out<=104;
				end
				if(in == 3) begin
					state<=5421;
					out<=105;
				end
				if(in == 4) begin
					state<=1532;
					out<=106;
				end
			end
			7343: begin
				if(in == 0) begin
					state<=7354;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=3465;
					out<=109;
				end
				if(in == 3) begin
					state<=5422;
					out<=110;
				end
				if(in == 4) begin
					state<=1533;
					out<=111;
				end
			end
			7344: begin
				if(in == 0) begin
					state<=7355;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=3466;
					out<=114;
				end
				if(in == 3) begin
					state<=5423;
					out<=115;
				end
				if(in == 4) begin
					state<=1534;
					out<=116;
				end
			end
			7345: begin
				if(in == 0) begin
					state<=7346;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=3457;
					out<=119;
				end
				if(in == 3) begin
					state<=5414;
					out<=120;
				end
				if(in == 4) begin
					state<=1525;
					out<=121;
				end
			end
			7346: begin
				if(in == 0) begin
					state<=7357;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=3468;
					out<=124;
				end
				if(in == 3) begin
					state<=5425;
					out<=125;
				end
				if(in == 4) begin
					state<=1536;
					out<=126;
				end
			end
			7347: begin
				if(in == 0) begin
					state<=7358;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=3469;
					out<=129;
				end
				if(in == 3) begin
					state<=5426;
					out<=130;
				end
				if(in == 4) begin
					state<=1537;
					out<=131;
				end
			end
			7348: begin
				if(in == 0) begin
					state<=7359;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=3470;
					out<=134;
				end
				if(in == 3) begin
					state<=5427;
					out<=135;
				end
				if(in == 4) begin
					state<=1538;
					out<=136;
				end
			end
			7349: begin
				if(in == 0) begin
					state<=7360;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=3471;
					out<=139;
				end
				if(in == 3) begin
					state<=5428;
					out<=140;
				end
				if(in == 4) begin
					state<=1539;
					out<=141;
				end
			end
			7350: begin
				if(in == 0) begin
					state<=7361;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=3472;
					out<=144;
				end
				if(in == 3) begin
					state<=5429;
					out<=145;
				end
				if(in == 4) begin
					state<=1540;
					out<=146;
				end
			end
			7351: begin
				if(in == 0) begin
					state<=7362;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=3473;
					out<=149;
				end
				if(in == 3) begin
					state<=5430;
					out<=150;
				end
				if(in == 4) begin
					state<=1541;
					out<=151;
				end
			end
			7352: begin
				if(in == 0) begin
					state<=7363;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=3474;
					out<=154;
				end
				if(in == 3) begin
					state<=5431;
					out<=155;
				end
				if(in == 4) begin
					state<=1542;
					out<=156;
				end
			end
			7353: begin
				if(in == 0) begin
					state<=7364;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=3475;
					out<=159;
				end
				if(in == 3) begin
					state<=5432;
					out<=160;
				end
				if(in == 4) begin
					state<=1543;
					out<=161;
				end
			end
			7354: begin
				if(in == 0) begin
					state<=7365;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=3476;
					out<=164;
				end
				if(in == 3) begin
					state<=5433;
					out<=165;
				end
				if(in == 4) begin
					state<=1544;
					out<=166;
				end
			end
			7355: begin
				if(in == 0) begin
					state<=7356;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=3467;
					out<=169;
				end
				if(in == 3) begin
					state<=5424;
					out<=170;
				end
				if(in == 4) begin
					state<=1535;
					out<=171;
				end
			end
			7356: begin
				if(in == 0) begin
					state<=6421;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=2532;
					out<=174;
				end
				if(in == 3) begin
					state<=4432;
					out<=175;
				end
				if(in == 4) begin
					state<=534;
					out<=176;
				end
			end
			7357: begin
				if(in == 0) begin
					state<=6422;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=2533;
					out<=179;
				end
				if(in == 3) begin
					state<=4433;
					out<=180;
				end
				if(in == 4) begin
					state<=535;
					out<=181;
				end
			end
			7358: begin
				if(in == 0) begin
					state<=6423;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=2534;
					out<=184;
				end
				if(in == 3) begin
					state<=4434;
					out<=185;
				end
				if(in == 4) begin
					state<=536;
					out<=186;
				end
			end
			7359: begin
				if(in == 0) begin
					state<=6424;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=2535;
					out<=189;
				end
				if(in == 3) begin
					state<=4435;
					out<=190;
				end
				if(in == 4) begin
					state<=537;
					out<=191;
				end
			end
			7360: begin
				if(in == 0) begin
					state<=6425;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=2536;
					out<=194;
				end
				if(in == 3) begin
					state<=4436;
					out<=195;
				end
				if(in == 4) begin
					state<=538;
					out<=196;
				end
			end
			7361: begin
				if(in == 0) begin
					state<=6426;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=2537;
					out<=199;
				end
				if(in == 3) begin
					state<=4437;
					out<=200;
				end
				if(in == 4) begin
					state<=539;
					out<=201;
				end
			end
			7362: begin
				if(in == 0) begin
					state<=6427;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=2538;
					out<=204;
				end
				if(in == 3) begin
					state<=4438;
					out<=205;
				end
				if(in == 4) begin
					state<=540;
					out<=206;
				end
			end
			7363: begin
				if(in == 0) begin
					state<=6428;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=2539;
					out<=209;
				end
				if(in == 3) begin
					state<=4439;
					out<=210;
				end
				if(in == 4) begin
					state<=541;
					out<=211;
				end
			end
			7364: begin
				if(in == 0) begin
					state<=6429;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=2540;
					out<=214;
				end
				if(in == 3) begin
					state<=4440;
					out<=215;
				end
				if(in == 4) begin
					state<=542;
					out<=216;
				end
			end
			7365: begin
				if(in == 0) begin
					state<=7366;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=3477;
					out<=219;
				end
				if(in == 3) begin
					state<=5434;
					out<=220;
				end
				if(in == 4) begin
					state<=1545;
					out<=221;
				end
			end
			7366: begin
				if(in == 0) begin
					state<=6431;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=2542;
					out<=224;
				end
				if(in == 3) begin
					state<=4442;
					out<=225;
				end
				if(in == 4) begin
					state<=544;
					out<=226;
				end
			end
			7367: begin
				if(in == 0) begin
					state<=7378;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=3489;
					out<=229;
				end
				if(in == 3) begin
					state<=5446;
					out<=230;
				end
				if(in == 4) begin
					state<=1557;
					out<=231;
				end
			end
			7368: begin
				if(in == 0) begin
					state<=7379;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=3490;
					out<=234;
				end
				if(in == 3) begin
					state<=5447;
					out<=235;
				end
				if(in == 4) begin
					state<=1558;
					out<=236;
				end
			end
			7369: begin
				if(in == 0) begin
					state<=7380;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=3491;
					out<=239;
				end
				if(in == 3) begin
					state<=5448;
					out<=240;
				end
				if(in == 4) begin
					state<=1559;
					out<=241;
				end
			end
			7370: begin
				if(in == 0) begin
					state<=7381;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=3492;
					out<=244;
				end
				if(in == 3) begin
					state<=5449;
					out<=245;
				end
				if(in == 4) begin
					state<=1560;
					out<=246;
				end
			end
			7371: begin
				if(in == 0) begin
					state<=7382;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=3493;
					out<=249;
				end
				if(in == 3) begin
					state<=5450;
					out<=250;
				end
				if(in == 4) begin
					state<=1561;
					out<=251;
				end
			end
			7372: begin
				if(in == 0) begin
					state<=7383;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=3494;
					out<=254;
				end
				if(in == 3) begin
					state<=5451;
					out<=255;
				end
				if(in == 4) begin
					state<=1562;
					out<=0;
				end
			end
			7373: begin
				if(in == 0) begin
					state<=7384;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=3495;
					out<=3;
				end
				if(in == 3) begin
					state<=5452;
					out<=4;
				end
				if(in == 4) begin
					state<=1563;
					out<=5;
				end
			end
			7374: begin
				if(in == 0) begin
					state<=7385;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=3496;
					out<=8;
				end
				if(in == 3) begin
					state<=5453;
					out<=9;
				end
				if(in == 4) begin
					state<=1564;
					out<=10;
				end
			end
			7375: begin
				if(in == 0) begin
					state<=7386;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=3497;
					out<=13;
				end
				if(in == 3) begin
					state<=5454;
					out<=14;
				end
				if(in == 4) begin
					state<=1565;
					out<=15;
				end
			end
			7376: begin
				if(in == 0) begin
					state<=7377;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=3488;
					out<=18;
				end
				if(in == 3) begin
					state<=5445;
					out<=19;
				end
				if(in == 4) begin
					state<=1556;
					out<=20;
				end
			end
			7377: begin
				if(in == 0) begin
					state<=7388;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=3499;
					out<=23;
				end
				if(in == 3) begin
					state<=5456;
					out<=24;
				end
				if(in == 4) begin
					state<=1567;
					out<=25;
				end
			end
			7378: begin
				if(in == 0) begin
					state<=7389;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=3500;
					out<=28;
				end
				if(in == 3) begin
					state<=5457;
					out<=29;
				end
				if(in == 4) begin
					state<=1568;
					out<=30;
				end
			end
			7379: begin
				if(in == 0) begin
					state<=7390;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=3501;
					out<=33;
				end
				if(in == 3) begin
					state<=5458;
					out<=34;
				end
				if(in == 4) begin
					state<=1569;
					out<=35;
				end
			end
			7380: begin
				if(in == 0) begin
					state<=7391;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=3502;
					out<=38;
				end
				if(in == 3) begin
					state<=5459;
					out<=39;
				end
				if(in == 4) begin
					state<=1570;
					out<=40;
				end
			end
			7381: begin
				if(in == 0) begin
					state<=7392;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=3503;
					out<=43;
				end
				if(in == 3) begin
					state<=5460;
					out<=44;
				end
				if(in == 4) begin
					state<=1571;
					out<=45;
				end
			end
			7382: begin
				if(in == 0) begin
					state<=7393;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=3504;
					out<=48;
				end
				if(in == 3) begin
					state<=5461;
					out<=49;
				end
				if(in == 4) begin
					state<=1572;
					out<=50;
				end
			end
			7383: begin
				if(in == 0) begin
					state<=7394;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=3505;
					out<=53;
				end
				if(in == 3) begin
					state<=5462;
					out<=54;
				end
				if(in == 4) begin
					state<=1573;
					out<=55;
				end
			end
			7384: begin
				if(in == 0) begin
					state<=7395;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=3506;
					out<=58;
				end
				if(in == 3) begin
					state<=5463;
					out<=59;
				end
				if(in == 4) begin
					state<=1574;
					out<=60;
				end
			end
			7385: begin
				if(in == 0) begin
					state<=7396;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=3507;
					out<=63;
				end
				if(in == 3) begin
					state<=5464;
					out<=64;
				end
				if(in == 4) begin
					state<=1575;
					out<=65;
				end
			end
			7386: begin
				if(in == 0) begin
					state<=7387;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=3498;
					out<=68;
				end
				if(in == 3) begin
					state<=5455;
					out<=69;
				end
				if(in == 4) begin
					state<=1566;
					out<=70;
				end
			end
			7387: begin
				if(in == 0) begin
					state<=6490;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=2601;
					out<=73;
				end
				if(in == 3) begin
					state<=4501;
					out<=74;
				end
				if(in == 4) begin
					state<=603;
					out<=75;
				end
			end
			7388: begin
				if(in == 0) begin
					state<=6491;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=2602;
					out<=78;
				end
				if(in == 3) begin
					state<=4502;
					out<=79;
				end
				if(in == 4) begin
					state<=604;
					out<=80;
				end
			end
			7389: begin
				if(in == 0) begin
					state<=6492;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=2603;
					out<=83;
				end
				if(in == 3) begin
					state<=4503;
					out<=84;
				end
				if(in == 4) begin
					state<=605;
					out<=85;
				end
			end
			7390: begin
				if(in == 0) begin
					state<=6493;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=2604;
					out<=88;
				end
				if(in == 3) begin
					state<=4504;
					out<=89;
				end
				if(in == 4) begin
					state<=606;
					out<=90;
				end
			end
			7391: begin
				if(in == 0) begin
					state<=6494;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=2605;
					out<=93;
				end
				if(in == 3) begin
					state<=4505;
					out<=94;
				end
				if(in == 4) begin
					state<=607;
					out<=95;
				end
			end
			7392: begin
				if(in == 0) begin
					state<=6495;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=2606;
					out<=98;
				end
				if(in == 3) begin
					state<=4506;
					out<=99;
				end
				if(in == 4) begin
					state<=608;
					out<=100;
				end
			end
			7393: begin
				if(in == 0) begin
					state<=6496;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=2607;
					out<=103;
				end
				if(in == 3) begin
					state<=4507;
					out<=104;
				end
				if(in == 4) begin
					state<=609;
					out<=105;
				end
			end
			7394: begin
				if(in == 0) begin
					state<=6497;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=2608;
					out<=108;
				end
				if(in == 3) begin
					state<=4508;
					out<=109;
				end
				if(in == 4) begin
					state<=610;
					out<=110;
				end
			end
			7395: begin
				if(in == 0) begin
					state<=6498;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=2609;
					out<=113;
				end
				if(in == 3) begin
					state<=4509;
					out<=114;
				end
				if(in == 4) begin
					state<=611;
					out<=115;
				end
			end
			7396: begin
				if(in == 0) begin
					state<=7397;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=3508;
					out<=118;
				end
				if(in == 3) begin
					state<=5465;
					out<=119;
				end
				if(in == 4) begin
					state<=1576;
					out<=120;
				end
			end
			7397: begin
				if(in == 0) begin
					state<=6500;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=2611;
					out<=123;
				end
				if(in == 3) begin
					state<=4511;
					out<=124;
				end
				if(in == 4) begin
					state<=613;
					out<=125;
				end
			end
			7398: begin
				if(in == 0) begin
					state<=7409;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=3520;
					out<=128;
				end
				if(in == 3) begin
					state<=5508;
					out<=129;
				end
				if(in == 4) begin
					state<=1619;
					out<=130;
				end
			end
			7399: begin
				if(in == 0) begin
					state<=7410;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=3521;
					out<=133;
				end
				if(in == 3) begin
					state<=5509;
					out<=134;
				end
				if(in == 4) begin
					state<=1620;
					out<=135;
				end
			end
			7400: begin
				if(in == 0) begin
					state<=7411;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=3522;
					out<=138;
				end
				if(in == 3) begin
					state<=5510;
					out<=139;
				end
				if(in == 4) begin
					state<=1621;
					out<=140;
				end
			end
			7401: begin
				if(in == 0) begin
					state<=7412;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=3523;
					out<=143;
				end
				if(in == 3) begin
					state<=5511;
					out<=144;
				end
				if(in == 4) begin
					state<=1622;
					out<=145;
				end
			end
			7402: begin
				if(in == 0) begin
					state<=7413;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=3524;
					out<=148;
				end
				if(in == 3) begin
					state<=5512;
					out<=149;
				end
				if(in == 4) begin
					state<=1623;
					out<=150;
				end
			end
			7403: begin
				if(in == 0) begin
					state<=7414;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=3525;
					out<=153;
				end
				if(in == 3) begin
					state<=5513;
					out<=154;
				end
				if(in == 4) begin
					state<=1624;
					out<=155;
				end
			end
			7404: begin
				if(in == 0) begin
					state<=7415;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=3526;
					out<=158;
				end
				if(in == 3) begin
					state<=5514;
					out<=159;
				end
				if(in == 4) begin
					state<=1625;
					out<=160;
				end
			end
			7405: begin
				if(in == 0) begin
					state<=7416;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=3527;
					out<=163;
				end
				if(in == 3) begin
					state<=5515;
					out<=164;
				end
				if(in == 4) begin
					state<=1626;
					out<=165;
				end
			end
			7406: begin
				if(in == 0) begin
					state<=7417;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=3528;
					out<=168;
				end
				if(in == 3) begin
					state<=5516;
					out<=169;
				end
				if(in == 4) begin
					state<=1627;
					out<=170;
				end
			end
			7407: begin
				if(in == 0) begin
					state<=7408;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=3519;
					out<=173;
				end
				if(in == 3) begin
					state<=5507;
					out<=174;
				end
				if(in == 4) begin
					state<=1618;
					out<=175;
				end
			end
			7408: begin
				if(in == 0) begin
					state<=7419;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=3530;
					out<=178;
				end
				if(in == 3) begin
					state<=5518;
					out<=179;
				end
				if(in == 4) begin
					state<=1629;
					out<=180;
				end
			end
			7409: begin
				if(in == 0) begin
					state<=7420;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=3531;
					out<=183;
				end
				if(in == 3) begin
					state<=5519;
					out<=184;
				end
				if(in == 4) begin
					state<=1630;
					out<=185;
				end
			end
			7410: begin
				if(in == 0) begin
					state<=7421;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=3532;
					out<=188;
				end
				if(in == 3) begin
					state<=5520;
					out<=189;
				end
				if(in == 4) begin
					state<=1631;
					out<=190;
				end
			end
			7411: begin
				if(in == 0) begin
					state<=7422;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=3533;
					out<=193;
				end
				if(in == 3) begin
					state<=5521;
					out<=194;
				end
				if(in == 4) begin
					state<=1632;
					out<=195;
				end
			end
			7412: begin
				if(in == 0) begin
					state<=7423;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=3534;
					out<=198;
				end
				if(in == 3) begin
					state<=5522;
					out<=199;
				end
				if(in == 4) begin
					state<=1633;
					out<=200;
				end
			end
			7413: begin
				if(in == 0) begin
					state<=7424;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=3535;
					out<=203;
				end
				if(in == 3) begin
					state<=5523;
					out<=204;
				end
				if(in == 4) begin
					state<=1634;
					out<=205;
				end
			end
			7414: begin
				if(in == 0) begin
					state<=7425;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=3536;
					out<=208;
				end
				if(in == 3) begin
					state<=5524;
					out<=209;
				end
				if(in == 4) begin
					state<=1635;
					out<=210;
				end
			end
			7415: begin
				if(in == 0) begin
					state<=7426;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=3537;
					out<=213;
				end
				if(in == 3) begin
					state<=5525;
					out<=214;
				end
				if(in == 4) begin
					state<=1636;
					out<=215;
				end
			end
			7416: begin
				if(in == 0) begin
					state<=7427;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=3538;
					out<=218;
				end
				if(in == 3) begin
					state<=5526;
					out<=219;
				end
				if(in == 4) begin
					state<=1637;
					out<=220;
				end
			end
			7417: begin
				if(in == 0) begin
					state<=7418;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=3529;
					out<=223;
				end
				if(in == 3) begin
					state<=5517;
					out<=224;
				end
				if(in == 4) begin
					state<=1628;
					out<=225;
				end
			end
			7418: begin
				if(in == 0) begin
					state<=7429;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=3540;
					out<=228;
				end
				if(in == 3) begin
					state<=5528;
					out<=229;
				end
				if(in == 4) begin
					state<=1639;
					out<=230;
				end
			end
			7419: begin
				if(in == 0) begin
					state<=7430;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=3541;
					out<=233;
				end
				if(in == 3) begin
					state<=5529;
					out<=234;
				end
				if(in == 4) begin
					state<=1640;
					out<=235;
				end
			end
			7420: begin
				if(in == 0) begin
					state<=7431;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=3542;
					out<=238;
				end
				if(in == 3) begin
					state<=5530;
					out<=239;
				end
				if(in == 4) begin
					state<=1641;
					out<=240;
				end
			end
			7421: begin
				if(in == 0) begin
					state<=7432;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=3543;
					out<=243;
				end
				if(in == 3) begin
					state<=5531;
					out<=244;
				end
				if(in == 4) begin
					state<=1642;
					out<=245;
				end
			end
			7422: begin
				if(in == 0) begin
					state<=7433;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=3544;
					out<=248;
				end
				if(in == 3) begin
					state<=5532;
					out<=249;
				end
				if(in == 4) begin
					state<=1643;
					out<=250;
				end
			end
			7423: begin
				if(in == 0) begin
					state<=7434;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=3545;
					out<=253;
				end
				if(in == 3) begin
					state<=5533;
					out<=254;
				end
				if(in == 4) begin
					state<=1644;
					out<=255;
				end
			end
			7424: begin
				if(in == 0) begin
					state<=7435;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=3546;
					out<=2;
				end
				if(in == 3) begin
					state<=5534;
					out<=3;
				end
				if(in == 4) begin
					state<=1645;
					out<=4;
				end
			end
			7425: begin
				if(in == 0) begin
					state<=7436;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=3547;
					out<=7;
				end
				if(in == 3) begin
					state<=5535;
					out<=8;
				end
				if(in == 4) begin
					state<=1646;
					out<=9;
				end
			end
			7426: begin
				if(in == 0) begin
					state<=7437;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=3548;
					out<=12;
				end
				if(in == 3) begin
					state<=5536;
					out<=13;
				end
				if(in == 4) begin
					state<=1647;
					out<=14;
				end
			end
			7427: begin
				if(in == 0) begin
					state<=7428;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=3539;
					out<=17;
				end
				if(in == 3) begin
					state<=5527;
					out<=18;
				end
				if(in == 4) begin
					state<=1638;
					out<=19;
				end
			end
			7428: begin
				if(in == 0) begin
					state<=7439;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=3550;
					out<=22;
				end
				if(in == 3) begin
					state<=5538;
					out<=23;
				end
				if(in == 4) begin
					state<=1649;
					out<=24;
				end
			end
			7429: begin
				if(in == 0) begin
					state<=7440;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=3551;
					out<=27;
				end
				if(in == 3) begin
					state<=5539;
					out<=28;
				end
				if(in == 4) begin
					state<=1650;
					out<=29;
				end
			end
			7430: begin
				if(in == 0) begin
					state<=7441;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=3552;
					out<=32;
				end
				if(in == 3) begin
					state<=5540;
					out<=33;
				end
				if(in == 4) begin
					state<=1651;
					out<=34;
				end
			end
			7431: begin
				if(in == 0) begin
					state<=7442;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=3553;
					out<=37;
				end
				if(in == 3) begin
					state<=5541;
					out<=38;
				end
				if(in == 4) begin
					state<=1652;
					out<=39;
				end
			end
			7432: begin
				if(in == 0) begin
					state<=7443;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=3554;
					out<=42;
				end
				if(in == 3) begin
					state<=5542;
					out<=43;
				end
				if(in == 4) begin
					state<=1653;
					out<=44;
				end
			end
			7433: begin
				if(in == 0) begin
					state<=7444;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=3555;
					out<=47;
				end
				if(in == 3) begin
					state<=5543;
					out<=48;
				end
				if(in == 4) begin
					state<=1654;
					out<=49;
				end
			end
			7434: begin
				if(in == 0) begin
					state<=7445;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=3556;
					out<=52;
				end
				if(in == 3) begin
					state<=5544;
					out<=53;
				end
				if(in == 4) begin
					state<=1655;
					out<=54;
				end
			end
			7435: begin
				if(in == 0) begin
					state<=7446;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=3557;
					out<=57;
				end
				if(in == 3) begin
					state<=5545;
					out<=58;
				end
				if(in == 4) begin
					state<=1656;
					out<=59;
				end
			end
			7436: begin
				if(in == 0) begin
					state<=7447;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=3558;
					out<=62;
				end
				if(in == 3) begin
					state<=5546;
					out<=63;
				end
				if(in == 4) begin
					state<=1657;
					out<=64;
				end
			end
			7437: begin
				if(in == 0) begin
					state<=7438;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=3549;
					out<=67;
				end
				if(in == 3) begin
					state<=5537;
					out<=68;
				end
				if(in == 4) begin
					state<=1648;
					out<=69;
				end
			end
			7438: begin
				if(in == 0) begin
					state<=7449;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=3560;
					out<=72;
				end
				if(in == 3) begin
					state<=5548;
					out<=73;
				end
				if(in == 4) begin
					state<=1659;
					out<=74;
				end
			end
			7439: begin
				if(in == 0) begin
					state<=7450;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=3561;
					out<=77;
				end
				if(in == 3) begin
					state<=5549;
					out<=78;
				end
				if(in == 4) begin
					state<=1660;
					out<=79;
				end
			end
			7440: begin
				if(in == 0) begin
					state<=7451;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=3562;
					out<=82;
				end
				if(in == 3) begin
					state<=5550;
					out<=83;
				end
				if(in == 4) begin
					state<=1661;
					out<=84;
				end
			end
			7441: begin
				if(in == 0) begin
					state<=7452;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=3563;
					out<=87;
				end
				if(in == 3) begin
					state<=5551;
					out<=88;
				end
				if(in == 4) begin
					state<=1662;
					out<=89;
				end
			end
			7442: begin
				if(in == 0) begin
					state<=7453;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=3564;
					out<=92;
				end
				if(in == 3) begin
					state<=5552;
					out<=93;
				end
				if(in == 4) begin
					state<=1663;
					out<=94;
				end
			end
			7443: begin
				if(in == 0) begin
					state<=7454;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=3565;
					out<=97;
				end
				if(in == 3) begin
					state<=5553;
					out<=98;
				end
				if(in == 4) begin
					state<=1664;
					out<=99;
				end
			end
			7444: begin
				if(in == 0) begin
					state<=7455;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=3566;
					out<=102;
				end
				if(in == 3) begin
					state<=5554;
					out<=103;
				end
				if(in == 4) begin
					state<=1665;
					out<=104;
				end
			end
			7445: begin
				if(in == 0) begin
					state<=7456;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=3567;
					out<=107;
				end
				if(in == 3) begin
					state<=5555;
					out<=108;
				end
				if(in == 4) begin
					state<=1666;
					out<=109;
				end
			end
			7446: begin
				if(in == 0) begin
					state<=7457;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=3568;
					out<=112;
				end
				if(in == 3) begin
					state<=5556;
					out<=113;
				end
				if(in == 4) begin
					state<=1667;
					out<=114;
				end
			end
			7447: begin
				if(in == 0) begin
					state<=7448;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=3559;
					out<=117;
				end
				if(in == 3) begin
					state<=5547;
					out<=118;
				end
				if(in == 4) begin
					state<=1658;
					out<=119;
				end
			end
			7448: begin
				if(in == 0) begin
					state<=7459;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=3570;
					out<=122;
				end
				if(in == 3) begin
					state<=5558;
					out<=123;
				end
				if(in == 4) begin
					state<=1669;
					out<=124;
				end
			end
			7449: begin
				if(in == 0) begin
					state<=7460;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=3571;
					out<=127;
				end
				if(in == 3) begin
					state<=5559;
					out<=128;
				end
				if(in == 4) begin
					state<=1670;
					out<=129;
				end
			end
			7450: begin
				if(in == 0) begin
					state<=7461;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=3572;
					out<=132;
				end
				if(in == 3) begin
					state<=5560;
					out<=133;
				end
				if(in == 4) begin
					state<=1671;
					out<=134;
				end
			end
			7451: begin
				if(in == 0) begin
					state<=7462;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=3573;
					out<=137;
				end
				if(in == 3) begin
					state<=5561;
					out<=138;
				end
				if(in == 4) begin
					state<=1672;
					out<=139;
				end
			end
			7452: begin
				if(in == 0) begin
					state<=7463;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=3574;
					out<=142;
				end
				if(in == 3) begin
					state<=5562;
					out<=143;
				end
				if(in == 4) begin
					state<=1673;
					out<=144;
				end
			end
			7453: begin
				if(in == 0) begin
					state<=7464;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=3575;
					out<=147;
				end
				if(in == 3) begin
					state<=5563;
					out<=148;
				end
				if(in == 4) begin
					state<=1674;
					out<=149;
				end
			end
			7454: begin
				if(in == 0) begin
					state<=7465;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=3576;
					out<=152;
				end
				if(in == 3) begin
					state<=5564;
					out<=153;
				end
				if(in == 4) begin
					state<=1675;
					out<=154;
				end
			end
			7455: begin
				if(in == 0) begin
					state<=7466;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=3577;
					out<=157;
				end
				if(in == 3) begin
					state<=5565;
					out<=158;
				end
				if(in == 4) begin
					state<=1676;
					out<=159;
				end
			end
			7456: begin
				if(in == 0) begin
					state<=7467;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=3578;
					out<=162;
				end
				if(in == 3) begin
					state<=5566;
					out<=163;
				end
				if(in == 4) begin
					state<=1677;
					out<=164;
				end
			end
			7457: begin
				if(in == 0) begin
					state<=7458;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=3569;
					out<=167;
				end
				if(in == 3) begin
					state<=5557;
					out<=168;
				end
				if(in == 4) begin
					state<=1668;
					out<=169;
				end
			end
			7458: begin
				if(in == 0) begin
					state<=7469;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=3580;
					out<=172;
				end
				if(in == 3) begin
					state<=5568;
					out<=173;
				end
				if(in == 4) begin
					state<=1679;
					out<=174;
				end
			end
			7459: begin
				if(in == 0) begin
					state<=7470;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=3581;
					out<=177;
				end
				if(in == 3) begin
					state<=5569;
					out<=178;
				end
				if(in == 4) begin
					state<=1680;
					out<=179;
				end
			end
			7460: begin
				if(in == 0) begin
					state<=7471;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=3582;
					out<=182;
				end
				if(in == 3) begin
					state<=5570;
					out<=183;
				end
				if(in == 4) begin
					state<=1681;
					out<=184;
				end
			end
			7461: begin
				if(in == 0) begin
					state<=7472;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=3583;
					out<=187;
				end
				if(in == 3) begin
					state<=5571;
					out<=188;
				end
				if(in == 4) begin
					state<=1682;
					out<=189;
				end
			end
			7462: begin
				if(in == 0) begin
					state<=7473;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=3584;
					out<=192;
				end
				if(in == 3) begin
					state<=5572;
					out<=193;
				end
				if(in == 4) begin
					state<=1683;
					out<=194;
				end
			end
			7463: begin
				if(in == 0) begin
					state<=7474;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=3585;
					out<=197;
				end
				if(in == 3) begin
					state<=5573;
					out<=198;
				end
				if(in == 4) begin
					state<=1684;
					out<=199;
				end
			end
			7464: begin
				if(in == 0) begin
					state<=7475;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=3586;
					out<=202;
				end
				if(in == 3) begin
					state<=5574;
					out<=203;
				end
				if(in == 4) begin
					state<=1685;
					out<=204;
				end
			end
			7465: begin
				if(in == 0) begin
					state<=7476;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=3587;
					out<=207;
				end
				if(in == 3) begin
					state<=5575;
					out<=208;
				end
				if(in == 4) begin
					state<=1686;
					out<=209;
				end
			end
			7466: begin
				if(in == 0) begin
					state<=7477;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=3588;
					out<=212;
				end
				if(in == 3) begin
					state<=5576;
					out<=213;
				end
				if(in == 4) begin
					state<=1687;
					out<=214;
				end
			end
			7467: begin
				if(in == 0) begin
					state<=7468;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=3579;
					out<=217;
				end
				if(in == 3) begin
					state<=5567;
					out<=218;
				end
				if(in == 4) begin
					state<=1678;
					out<=219;
				end
			end
			7468: begin
				if(in == 0) begin
					state<=7479;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=3590;
					out<=222;
				end
				if(in == 3) begin
					state<=5578;
					out<=223;
				end
				if(in == 4) begin
					state<=1689;
					out<=224;
				end
			end
			7469: begin
				if(in == 0) begin
					state<=7480;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=3591;
					out<=227;
				end
				if(in == 3) begin
					state<=5579;
					out<=228;
				end
				if(in == 4) begin
					state<=1690;
					out<=229;
				end
			end
			7470: begin
				if(in == 0) begin
					state<=7481;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=3592;
					out<=232;
				end
				if(in == 3) begin
					state<=5580;
					out<=233;
				end
				if(in == 4) begin
					state<=1691;
					out<=234;
				end
			end
			7471: begin
				if(in == 0) begin
					state<=7482;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=3593;
					out<=237;
				end
				if(in == 3) begin
					state<=5581;
					out<=238;
				end
				if(in == 4) begin
					state<=1692;
					out<=239;
				end
			end
			7472: begin
				if(in == 0) begin
					state<=7483;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=3594;
					out<=242;
				end
				if(in == 3) begin
					state<=5582;
					out<=243;
				end
				if(in == 4) begin
					state<=1693;
					out<=244;
				end
			end
			7473: begin
				if(in == 0) begin
					state<=7484;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=3595;
					out<=247;
				end
				if(in == 3) begin
					state<=5583;
					out<=248;
				end
				if(in == 4) begin
					state<=1694;
					out<=249;
				end
			end
			7474: begin
				if(in == 0) begin
					state<=7485;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=3596;
					out<=252;
				end
				if(in == 3) begin
					state<=5584;
					out<=253;
				end
				if(in == 4) begin
					state<=1695;
					out<=254;
				end
			end
			7475: begin
				if(in == 0) begin
					state<=7486;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=3597;
					out<=1;
				end
				if(in == 3) begin
					state<=5585;
					out<=2;
				end
				if(in == 4) begin
					state<=1696;
					out<=3;
				end
			end
			7476: begin
				if(in == 0) begin
					state<=7487;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=3598;
					out<=6;
				end
				if(in == 3) begin
					state<=5586;
					out<=7;
				end
				if(in == 4) begin
					state<=1697;
					out<=8;
				end
			end
			7477: begin
				if(in == 0) begin
					state<=7478;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=3589;
					out<=11;
				end
				if(in == 3) begin
					state<=5577;
					out<=12;
				end
				if(in == 4) begin
					state<=1688;
					out<=13;
				end
			end
			7478: begin
				if(in == 0) begin
					state<=7489;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=3600;
					out<=16;
				end
				if(in == 3) begin
					state<=5588;
					out<=17;
				end
				if(in == 4) begin
					state<=1699;
					out<=18;
				end
			end
			7479: begin
				if(in == 0) begin
					state<=7490;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=3601;
					out<=21;
				end
				if(in == 3) begin
					state<=5589;
					out<=22;
				end
				if(in == 4) begin
					state<=1700;
					out<=23;
				end
			end
			7480: begin
				if(in == 0) begin
					state<=7491;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=3602;
					out<=26;
				end
				if(in == 3) begin
					state<=5590;
					out<=27;
				end
				if(in == 4) begin
					state<=1701;
					out<=28;
				end
			end
			7481: begin
				if(in == 0) begin
					state<=7492;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=3603;
					out<=31;
				end
				if(in == 3) begin
					state<=5591;
					out<=32;
				end
				if(in == 4) begin
					state<=1702;
					out<=33;
				end
			end
			7482: begin
				if(in == 0) begin
					state<=7493;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=3604;
					out<=36;
				end
				if(in == 3) begin
					state<=5592;
					out<=37;
				end
				if(in == 4) begin
					state<=1703;
					out<=38;
				end
			end
			7483: begin
				if(in == 0) begin
					state<=7494;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=3605;
					out<=41;
				end
				if(in == 3) begin
					state<=5593;
					out<=42;
				end
				if(in == 4) begin
					state<=1704;
					out<=43;
				end
			end
			7484: begin
				if(in == 0) begin
					state<=7495;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=3606;
					out<=46;
				end
				if(in == 3) begin
					state<=5594;
					out<=47;
				end
				if(in == 4) begin
					state<=1705;
					out<=48;
				end
			end
			7485: begin
				if(in == 0) begin
					state<=7496;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=3607;
					out<=51;
				end
				if(in == 3) begin
					state<=5595;
					out<=52;
				end
				if(in == 4) begin
					state<=1706;
					out<=53;
				end
			end
			7486: begin
				if(in == 0) begin
					state<=7497;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=3608;
					out<=56;
				end
				if(in == 3) begin
					state<=5596;
					out<=57;
				end
				if(in == 4) begin
					state<=1707;
					out<=58;
				end
			end
			7487: begin
				if(in == 0) begin
					state<=7488;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=3599;
					out<=61;
				end
				if(in == 3) begin
					state<=5587;
					out<=62;
				end
				if(in == 4) begin
					state<=1698;
					out<=63;
				end
			end
			7488: begin
				if(in == 0) begin
					state<=7499;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=3610;
					out<=66;
				end
				if(in == 3) begin
					state<=5598;
					out<=67;
				end
				if(in == 4) begin
					state<=1709;
					out<=68;
				end
			end
			7489: begin
				if(in == 0) begin
					state<=7500;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=3611;
					out<=71;
				end
				if(in == 3) begin
					state<=5599;
					out<=72;
				end
				if(in == 4) begin
					state<=1710;
					out<=73;
				end
			end
			7490: begin
				if(in == 0) begin
					state<=7501;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=3612;
					out<=76;
				end
				if(in == 3) begin
					state<=5600;
					out<=77;
				end
				if(in == 4) begin
					state<=1711;
					out<=78;
				end
			end
			7491: begin
				if(in == 0) begin
					state<=7502;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=3613;
					out<=81;
				end
				if(in == 3) begin
					state<=5601;
					out<=82;
				end
				if(in == 4) begin
					state<=1712;
					out<=83;
				end
			end
			7492: begin
				if(in == 0) begin
					state<=7503;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=3614;
					out<=86;
				end
				if(in == 3) begin
					state<=5602;
					out<=87;
				end
				if(in == 4) begin
					state<=1713;
					out<=88;
				end
			end
			7493: begin
				if(in == 0) begin
					state<=7504;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=3615;
					out<=91;
				end
				if(in == 3) begin
					state<=5603;
					out<=92;
				end
				if(in == 4) begin
					state<=1714;
					out<=93;
				end
			end
			7494: begin
				if(in == 0) begin
					state<=7505;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=3616;
					out<=96;
				end
				if(in == 3) begin
					state<=5604;
					out<=97;
				end
				if(in == 4) begin
					state<=1715;
					out<=98;
				end
			end
			7495: begin
				if(in == 0) begin
					state<=7506;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=3617;
					out<=101;
				end
				if(in == 3) begin
					state<=5605;
					out<=102;
				end
				if(in == 4) begin
					state<=1716;
					out<=103;
				end
			end
			7496: begin
				if(in == 0) begin
					state<=7507;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=3618;
					out<=106;
				end
				if(in == 3) begin
					state<=5606;
					out<=107;
				end
				if(in == 4) begin
					state<=1717;
					out<=108;
				end
			end
			7497: begin
				if(in == 0) begin
					state<=7498;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=3609;
					out<=111;
				end
				if(in == 3) begin
					state<=5597;
					out<=112;
				end
				if(in == 4) begin
					state<=1708;
					out<=113;
				end
			end
			7498: begin
				if(in == 0) begin
					state<=7509;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=3620;
					out<=116;
				end
				if(in == 3) begin
					state<=5608;
					out<=117;
				end
				if(in == 4) begin
					state<=1719;
					out<=118;
				end
			end
			7499: begin
				if(in == 0) begin
					state<=7510;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=3621;
					out<=121;
				end
				if(in == 3) begin
					state<=5609;
					out<=122;
				end
				if(in == 4) begin
					state<=1720;
					out<=123;
				end
			end
			7500: begin
				if(in == 0) begin
					state<=7511;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=3622;
					out<=126;
				end
				if(in == 3) begin
					state<=5610;
					out<=127;
				end
				if(in == 4) begin
					state<=1721;
					out<=128;
				end
			end
			7501: begin
				if(in == 0) begin
					state<=7512;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=3623;
					out<=131;
				end
				if(in == 3) begin
					state<=5611;
					out<=132;
				end
				if(in == 4) begin
					state<=1722;
					out<=133;
				end
			end
			7502: begin
				if(in == 0) begin
					state<=7513;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=3624;
					out<=136;
				end
				if(in == 3) begin
					state<=5612;
					out<=137;
				end
				if(in == 4) begin
					state<=1723;
					out<=138;
				end
			end
			7503: begin
				if(in == 0) begin
					state<=7514;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=3625;
					out<=141;
				end
				if(in == 3) begin
					state<=5613;
					out<=142;
				end
				if(in == 4) begin
					state<=1724;
					out<=143;
				end
			end
			7504: begin
				if(in == 0) begin
					state<=7515;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=3626;
					out<=146;
				end
				if(in == 3) begin
					state<=5614;
					out<=147;
				end
				if(in == 4) begin
					state<=1725;
					out<=148;
				end
			end
			7505: begin
				if(in == 0) begin
					state<=7516;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=3627;
					out<=151;
				end
				if(in == 3) begin
					state<=5615;
					out<=152;
				end
				if(in == 4) begin
					state<=1726;
					out<=153;
				end
			end
			7506: begin
				if(in == 0) begin
					state<=7517;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=3628;
					out<=156;
				end
				if(in == 3) begin
					state<=5616;
					out<=157;
				end
				if(in == 4) begin
					state<=1727;
					out<=158;
				end
			end
			7507: begin
				if(in == 0) begin
					state<=7508;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=3619;
					out<=161;
				end
				if(in == 3) begin
					state<=5607;
					out<=162;
				end
				if(in == 4) begin
					state<=1718;
					out<=163;
				end
			end
			7508: begin
				if(in == 0) begin
					state<=7519;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=3630;
					out<=166;
				end
				if(in == 3) begin
					state<=5618;
					out<=167;
				end
				if(in == 4) begin
					state<=1729;
					out<=168;
				end
			end
			7509: begin
				if(in == 0) begin
					state<=7520;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=3631;
					out<=171;
				end
				if(in == 3) begin
					state<=5619;
					out<=172;
				end
				if(in == 4) begin
					state<=1730;
					out<=173;
				end
			end
			7510: begin
				if(in == 0) begin
					state<=7521;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=3632;
					out<=176;
				end
				if(in == 3) begin
					state<=5620;
					out<=177;
				end
				if(in == 4) begin
					state<=1731;
					out<=178;
				end
			end
			7511: begin
				if(in == 0) begin
					state<=7522;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=3633;
					out<=181;
				end
				if(in == 3) begin
					state<=5621;
					out<=182;
				end
				if(in == 4) begin
					state<=1732;
					out<=183;
				end
			end
			7512: begin
				if(in == 0) begin
					state<=7523;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=3634;
					out<=186;
				end
				if(in == 3) begin
					state<=5622;
					out<=187;
				end
				if(in == 4) begin
					state<=1733;
					out<=188;
				end
			end
			7513: begin
				if(in == 0) begin
					state<=7524;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=3635;
					out<=191;
				end
				if(in == 3) begin
					state<=5623;
					out<=192;
				end
				if(in == 4) begin
					state<=1734;
					out<=193;
				end
			end
			7514: begin
				if(in == 0) begin
					state<=7525;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=3636;
					out<=196;
				end
				if(in == 3) begin
					state<=5624;
					out<=197;
				end
				if(in == 4) begin
					state<=1735;
					out<=198;
				end
			end
			7515: begin
				if(in == 0) begin
					state<=7526;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=3637;
					out<=201;
				end
				if(in == 3) begin
					state<=5625;
					out<=202;
				end
				if(in == 4) begin
					state<=1736;
					out<=203;
				end
			end
			7516: begin
				if(in == 0) begin
					state<=7527;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=3638;
					out<=206;
				end
				if(in == 3) begin
					state<=5626;
					out<=207;
				end
				if(in == 4) begin
					state<=1737;
					out<=208;
				end
			end
			7517: begin
				if(in == 0) begin
					state<=7518;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=3629;
					out<=211;
				end
				if(in == 3) begin
					state<=5617;
					out<=212;
				end
				if(in == 4) begin
					state<=1728;
					out<=213;
				end
			end
			7518: begin
				if(in == 0) begin
					state<=7529;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=3640;
					out<=216;
				end
				if(in == 3) begin
					state<=5628;
					out<=217;
				end
				if(in == 4) begin
					state<=1739;
					out<=218;
				end
			end
			7519: begin
				if(in == 0) begin
					state<=7530;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=3641;
					out<=221;
				end
				if(in == 3) begin
					state<=5629;
					out<=222;
				end
				if(in == 4) begin
					state<=1740;
					out<=223;
				end
			end
			7520: begin
				if(in == 0) begin
					state<=7531;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=3642;
					out<=226;
				end
				if(in == 3) begin
					state<=5630;
					out<=227;
				end
				if(in == 4) begin
					state<=1741;
					out<=228;
				end
			end
			7521: begin
				if(in == 0) begin
					state<=7532;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=3643;
					out<=231;
				end
				if(in == 3) begin
					state<=5631;
					out<=232;
				end
				if(in == 4) begin
					state<=1742;
					out<=233;
				end
			end
			7522: begin
				if(in == 0) begin
					state<=7533;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=3644;
					out<=236;
				end
				if(in == 3) begin
					state<=5632;
					out<=237;
				end
				if(in == 4) begin
					state<=1743;
					out<=238;
				end
			end
			7523: begin
				if(in == 0) begin
					state<=7534;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=3645;
					out<=241;
				end
				if(in == 3) begin
					state<=5633;
					out<=242;
				end
				if(in == 4) begin
					state<=1744;
					out<=243;
				end
			end
			7524: begin
				if(in == 0) begin
					state<=7535;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=3646;
					out<=246;
				end
				if(in == 3) begin
					state<=5634;
					out<=247;
				end
				if(in == 4) begin
					state<=1745;
					out<=248;
				end
			end
			7525: begin
				if(in == 0) begin
					state<=7536;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=3647;
					out<=251;
				end
				if(in == 3) begin
					state<=5635;
					out<=252;
				end
				if(in == 4) begin
					state<=1746;
					out<=253;
				end
			end
			7526: begin
				if(in == 0) begin
					state<=7537;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=3648;
					out<=0;
				end
				if(in == 3) begin
					state<=5636;
					out<=1;
				end
				if(in == 4) begin
					state<=1747;
					out<=2;
				end
			end
			7527: begin
				if(in == 0) begin
					state<=7528;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=3639;
					out<=5;
				end
				if(in == 3) begin
					state<=5627;
					out<=6;
				end
				if(in == 4) begin
					state<=1738;
					out<=7;
				end
			end
			7528: begin
				if(in == 0) begin
					state<=7539;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=3650;
					out<=10;
				end
				if(in == 3) begin
					state<=5638;
					out<=11;
				end
				if(in == 4) begin
					state<=1749;
					out<=12;
				end
			end
			7529: begin
				if(in == 0) begin
					state<=7540;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=3651;
					out<=15;
				end
				if(in == 3) begin
					state<=5639;
					out<=16;
				end
				if(in == 4) begin
					state<=1750;
					out<=17;
				end
			end
			7530: begin
				if(in == 0) begin
					state<=7541;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=3652;
					out<=20;
				end
				if(in == 3) begin
					state<=5640;
					out<=21;
				end
				if(in == 4) begin
					state<=1751;
					out<=22;
				end
			end
			7531: begin
				if(in == 0) begin
					state<=7542;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=3653;
					out<=25;
				end
				if(in == 3) begin
					state<=5641;
					out<=26;
				end
				if(in == 4) begin
					state<=1752;
					out<=27;
				end
			end
			7532: begin
				if(in == 0) begin
					state<=7543;
					out<=28;
				end
				if(in == 1) begin
					state<=800;
					out<=29;
				end
				if(in == 2) begin
					state<=3654;
					out<=30;
				end
				if(in == 3) begin
					state<=5642;
					out<=31;
				end
				if(in == 4) begin
					state<=1753;
					out<=32;
				end
			end
			7533: begin
				if(in == 0) begin
					state<=7544;
					out<=33;
				end
				if(in == 1) begin
					state<=800;
					out<=34;
				end
				if(in == 2) begin
					state<=3655;
					out<=35;
				end
				if(in == 3) begin
					state<=5643;
					out<=36;
				end
				if(in == 4) begin
					state<=1754;
					out<=37;
				end
			end
			7534: begin
				if(in == 0) begin
					state<=7545;
					out<=38;
				end
				if(in == 1) begin
					state<=800;
					out<=39;
				end
				if(in == 2) begin
					state<=3656;
					out<=40;
				end
				if(in == 3) begin
					state<=5644;
					out<=41;
				end
				if(in == 4) begin
					state<=1755;
					out<=42;
				end
			end
			7535: begin
				if(in == 0) begin
					state<=7546;
					out<=43;
				end
				if(in == 1) begin
					state<=800;
					out<=44;
				end
				if(in == 2) begin
					state<=3657;
					out<=45;
				end
				if(in == 3) begin
					state<=5645;
					out<=46;
				end
				if(in == 4) begin
					state<=1756;
					out<=47;
				end
			end
			7536: begin
				if(in == 0) begin
					state<=7547;
					out<=48;
				end
				if(in == 1) begin
					state<=800;
					out<=49;
				end
				if(in == 2) begin
					state<=3658;
					out<=50;
				end
				if(in == 3) begin
					state<=5646;
					out<=51;
				end
				if(in == 4) begin
					state<=1757;
					out<=52;
				end
			end
			7537: begin
				if(in == 0) begin
					state<=7538;
					out<=53;
				end
				if(in == 1) begin
					state<=800;
					out<=54;
				end
				if(in == 2) begin
					state<=3649;
					out<=55;
				end
				if(in == 3) begin
					state<=5637;
					out<=56;
				end
				if(in == 4) begin
					state<=1748;
					out<=57;
				end
			end
			7538: begin
				if(in == 0) begin
					state<=7549;
					out<=58;
				end
				if(in == 1) begin
					state<=800;
					out<=59;
				end
				if(in == 2) begin
					state<=3660;
					out<=60;
				end
				if(in == 3) begin
					state<=5648;
					out<=61;
				end
				if(in == 4) begin
					state<=1759;
					out<=62;
				end
			end
			7539: begin
				if(in == 0) begin
					state<=7550;
					out<=63;
				end
				if(in == 1) begin
					state<=800;
					out<=64;
				end
				if(in == 2) begin
					state<=3661;
					out<=65;
				end
				if(in == 3) begin
					state<=5649;
					out<=66;
				end
				if(in == 4) begin
					state<=1760;
					out<=67;
				end
			end
			7540: begin
				if(in == 0) begin
					state<=7551;
					out<=68;
				end
				if(in == 1) begin
					state<=800;
					out<=69;
				end
				if(in == 2) begin
					state<=3662;
					out<=70;
				end
				if(in == 3) begin
					state<=5650;
					out<=71;
				end
				if(in == 4) begin
					state<=1761;
					out<=72;
				end
			end
			7541: begin
				if(in == 0) begin
					state<=7552;
					out<=73;
				end
				if(in == 1) begin
					state<=800;
					out<=74;
				end
				if(in == 2) begin
					state<=3663;
					out<=75;
				end
				if(in == 3) begin
					state<=5651;
					out<=76;
				end
				if(in == 4) begin
					state<=1762;
					out<=77;
				end
			end
			7542: begin
				if(in == 0) begin
					state<=7553;
					out<=78;
				end
				if(in == 1) begin
					state<=800;
					out<=79;
				end
				if(in == 2) begin
					state<=3664;
					out<=80;
				end
				if(in == 3) begin
					state<=5652;
					out<=81;
				end
				if(in == 4) begin
					state<=1763;
					out<=82;
				end
			end
			7543: begin
				if(in == 0) begin
					state<=7554;
					out<=83;
				end
				if(in == 1) begin
					state<=800;
					out<=84;
				end
				if(in == 2) begin
					state<=3665;
					out<=85;
				end
				if(in == 3) begin
					state<=5653;
					out<=86;
				end
				if(in == 4) begin
					state<=1764;
					out<=87;
				end
			end
			7544: begin
				if(in == 0) begin
					state<=7555;
					out<=88;
				end
				if(in == 1) begin
					state<=800;
					out<=89;
				end
				if(in == 2) begin
					state<=3666;
					out<=90;
				end
				if(in == 3) begin
					state<=5654;
					out<=91;
				end
				if(in == 4) begin
					state<=1765;
					out<=92;
				end
			end
			7545: begin
				if(in == 0) begin
					state<=7556;
					out<=93;
				end
				if(in == 1) begin
					state<=800;
					out<=94;
				end
				if(in == 2) begin
					state<=3667;
					out<=95;
				end
				if(in == 3) begin
					state<=5655;
					out<=96;
				end
				if(in == 4) begin
					state<=1766;
					out<=97;
				end
			end
			7546: begin
				if(in == 0) begin
					state<=7557;
					out<=98;
				end
				if(in == 1) begin
					state<=800;
					out<=99;
				end
				if(in == 2) begin
					state<=3668;
					out<=100;
				end
				if(in == 3) begin
					state<=5656;
					out<=101;
				end
				if(in == 4) begin
					state<=1767;
					out<=102;
				end
			end
			7547: begin
				if(in == 0) begin
					state<=7548;
					out<=103;
				end
				if(in == 1) begin
					state<=800;
					out<=104;
				end
				if(in == 2) begin
					state<=3659;
					out<=105;
				end
				if(in == 3) begin
					state<=5647;
					out<=106;
				end
				if(in == 4) begin
					state<=1758;
					out<=107;
				end
			end
			7548: begin
				if(in == 0) begin
					state<=7559;
					out<=108;
				end
				if(in == 1) begin
					state<=800;
					out<=109;
				end
				if(in == 2) begin
					state<=3670;
					out<=110;
				end
				if(in == 3) begin
					state<=5658;
					out<=111;
				end
				if(in == 4) begin
					state<=1769;
					out<=112;
				end
			end
			7549: begin
				if(in == 0) begin
					state<=7560;
					out<=113;
				end
				if(in == 1) begin
					state<=800;
					out<=114;
				end
				if(in == 2) begin
					state<=3671;
					out<=115;
				end
				if(in == 3) begin
					state<=5659;
					out<=116;
				end
				if(in == 4) begin
					state<=1770;
					out<=117;
				end
			end
			7550: begin
				if(in == 0) begin
					state<=7561;
					out<=118;
				end
				if(in == 1) begin
					state<=800;
					out<=119;
				end
				if(in == 2) begin
					state<=3672;
					out<=120;
				end
				if(in == 3) begin
					state<=5660;
					out<=121;
				end
				if(in == 4) begin
					state<=1771;
					out<=122;
				end
			end
			7551: begin
				if(in == 0) begin
					state<=7562;
					out<=123;
				end
				if(in == 1) begin
					state<=800;
					out<=124;
				end
				if(in == 2) begin
					state<=3673;
					out<=125;
				end
				if(in == 3) begin
					state<=5661;
					out<=126;
				end
				if(in == 4) begin
					state<=1772;
					out<=127;
				end
			end
			7552: begin
				if(in == 0) begin
					state<=7563;
					out<=128;
				end
				if(in == 1) begin
					state<=800;
					out<=129;
				end
				if(in == 2) begin
					state<=3674;
					out<=130;
				end
				if(in == 3) begin
					state<=5662;
					out<=131;
				end
				if(in == 4) begin
					state<=1773;
					out<=132;
				end
			end
			7553: begin
				if(in == 0) begin
					state<=7564;
					out<=133;
				end
				if(in == 1) begin
					state<=800;
					out<=134;
				end
				if(in == 2) begin
					state<=3675;
					out<=135;
				end
				if(in == 3) begin
					state<=5663;
					out<=136;
				end
				if(in == 4) begin
					state<=1774;
					out<=137;
				end
			end
			7554: begin
				if(in == 0) begin
					state<=7565;
					out<=138;
				end
				if(in == 1) begin
					state<=800;
					out<=139;
				end
				if(in == 2) begin
					state<=3676;
					out<=140;
				end
				if(in == 3) begin
					state<=5664;
					out<=141;
				end
				if(in == 4) begin
					state<=1775;
					out<=142;
				end
			end
			7555: begin
				if(in == 0) begin
					state<=7566;
					out<=143;
				end
				if(in == 1) begin
					state<=800;
					out<=144;
				end
				if(in == 2) begin
					state<=3677;
					out<=145;
				end
				if(in == 3) begin
					state<=5665;
					out<=146;
				end
				if(in == 4) begin
					state<=1776;
					out<=147;
				end
			end
			7556: begin
				if(in == 0) begin
					state<=7567;
					out<=148;
				end
				if(in == 1) begin
					state<=800;
					out<=149;
				end
				if(in == 2) begin
					state<=3678;
					out<=150;
				end
				if(in == 3) begin
					state<=5666;
					out<=151;
				end
				if(in == 4) begin
					state<=1777;
					out<=152;
				end
			end
			7557: begin
				if(in == 0) begin
					state<=7558;
					out<=153;
				end
				if(in == 1) begin
					state<=800;
					out<=154;
				end
				if(in == 2) begin
					state<=3669;
					out<=155;
				end
				if(in == 3) begin
					state<=5657;
					out<=156;
				end
				if(in == 4) begin
					state<=1768;
					out<=157;
				end
			end
			7558: begin
				if(in == 0) begin
					state<=7569;
					out<=158;
				end
				if(in == 1) begin
					state<=800;
					out<=159;
				end
				if(in == 2) begin
					state<=3680;
					out<=160;
				end
				if(in == 3) begin
					state<=5668;
					out<=161;
				end
				if(in == 4) begin
					state<=1779;
					out<=162;
				end
			end
			7559: begin
				if(in == 0) begin
					state<=7570;
					out<=163;
				end
				if(in == 1) begin
					state<=800;
					out<=164;
				end
				if(in == 2) begin
					state<=3681;
					out<=165;
				end
				if(in == 3) begin
					state<=5669;
					out<=166;
				end
				if(in == 4) begin
					state<=1780;
					out<=167;
				end
			end
			7560: begin
				if(in == 0) begin
					state<=7571;
					out<=168;
				end
				if(in == 1) begin
					state<=800;
					out<=169;
				end
				if(in == 2) begin
					state<=3682;
					out<=170;
				end
				if(in == 3) begin
					state<=5670;
					out<=171;
				end
				if(in == 4) begin
					state<=1781;
					out<=172;
				end
			end
			7561: begin
				if(in == 0) begin
					state<=7572;
					out<=173;
				end
				if(in == 1) begin
					state<=800;
					out<=174;
				end
				if(in == 2) begin
					state<=3683;
					out<=175;
				end
				if(in == 3) begin
					state<=5671;
					out<=176;
				end
				if(in == 4) begin
					state<=1782;
					out<=177;
				end
			end
			7562: begin
				if(in == 0) begin
					state<=7573;
					out<=178;
				end
				if(in == 1) begin
					state<=800;
					out<=179;
				end
				if(in == 2) begin
					state<=3684;
					out<=180;
				end
				if(in == 3) begin
					state<=5672;
					out<=181;
				end
				if(in == 4) begin
					state<=1783;
					out<=182;
				end
			end
			7563: begin
				if(in == 0) begin
					state<=7574;
					out<=183;
				end
				if(in == 1) begin
					state<=800;
					out<=184;
				end
				if(in == 2) begin
					state<=3685;
					out<=185;
				end
				if(in == 3) begin
					state<=5673;
					out<=186;
				end
				if(in == 4) begin
					state<=1784;
					out<=187;
				end
			end
			7564: begin
				if(in == 0) begin
					state<=7575;
					out<=188;
				end
				if(in == 1) begin
					state<=800;
					out<=189;
				end
				if(in == 2) begin
					state<=3686;
					out<=190;
				end
				if(in == 3) begin
					state<=5674;
					out<=191;
				end
				if(in == 4) begin
					state<=1785;
					out<=192;
				end
			end
			7565: begin
				if(in == 0) begin
					state<=7576;
					out<=193;
				end
				if(in == 1) begin
					state<=800;
					out<=194;
				end
				if(in == 2) begin
					state<=3687;
					out<=195;
				end
				if(in == 3) begin
					state<=5675;
					out<=196;
				end
				if(in == 4) begin
					state<=1786;
					out<=197;
				end
			end
			7566: begin
				if(in == 0) begin
					state<=7577;
					out<=198;
				end
				if(in == 1) begin
					state<=800;
					out<=199;
				end
				if(in == 2) begin
					state<=3688;
					out<=200;
				end
				if(in == 3) begin
					state<=5676;
					out<=201;
				end
				if(in == 4) begin
					state<=1787;
					out<=202;
				end
			end
			7567: begin
				if(in == 0) begin
					state<=7568;
					out<=203;
				end
				if(in == 1) begin
					state<=800;
					out<=204;
				end
				if(in == 2) begin
					state<=3679;
					out<=205;
				end
				if(in == 3) begin
					state<=5667;
					out<=206;
				end
				if(in == 4) begin
					state<=1778;
					out<=207;
				end
			end
			7568: begin
				if(in == 0) begin
					state<=7579;
					out<=208;
				end
				if(in == 1) begin
					state<=800;
					out<=209;
				end
				if(in == 2) begin
					state<=3690;
					out<=210;
				end
				if(in == 3) begin
					state<=5678;
					out<=211;
				end
				if(in == 4) begin
					state<=1789;
					out<=212;
				end
			end
			7569: begin
				if(in == 0) begin
					state<=7580;
					out<=213;
				end
				if(in == 1) begin
					state<=800;
					out<=214;
				end
				if(in == 2) begin
					state<=3691;
					out<=215;
				end
				if(in == 3) begin
					state<=5679;
					out<=216;
				end
				if(in == 4) begin
					state<=1790;
					out<=217;
				end
			end
			7570: begin
				if(in == 0) begin
					state<=7581;
					out<=218;
				end
				if(in == 1) begin
					state<=800;
					out<=219;
				end
				if(in == 2) begin
					state<=3692;
					out<=220;
				end
				if(in == 3) begin
					state<=5680;
					out<=221;
				end
				if(in == 4) begin
					state<=1791;
					out<=222;
				end
			end
			7571: begin
				if(in == 0) begin
					state<=7582;
					out<=223;
				end
				if(in == 1) begin
					state<=800;
					out<=224;
				end
				if(in == 2) begin
					state<=3693;
					out<=225;
				end
				if(in == 3) begin
					state<=5681;
					out<=226;
				end
				if(in == 4) begin
					state<=1792;
					out<=227;
				end
			end
			7572: begin
				if(in == 0) begin
					state<=7583;
					out<=228;
				end
				if(in == 1) begin
					state<=800;
					out<=229;
				end
				if(in == 2) begin
					state<=3694;
					out<=230;
				end
				if(in == 3) begin
					state<=5682;
					out<=231;
				end
				if(in == 4) begin
					state<=1793;
					out<=232;
				end
			end
			7573: begin
				if(in == 0) begin
					state<=7584;
					out<=233;
				end
				if(in == 1) begin
					state<=800;
					out<=234;
				end
				if(in == 2) begin
					state<=3695;
					out<=235;
				end
				if(in == 3) begin
					state<=5683;
					out<=236;
				end
				if(in == 4) begin
					state<=1794;
					out<=237;
				end
			end
			7574: begin
				if(in == 0) begin
					state<=7585;
					out<=238;
				end
				if(in == 1) begin
					state<=800;
					out<=239;
				end
				if(in == 2) begin
					state<=3696;
					out<=240;
				end
				if(in == 3) begin
					state<=5684;
					out<=241;
				end
				if(in == 4) begin
					state<=1795;
					out<=242;
				end
			end
			7575: begin
				if(in == 0) begin
					state<=7586;
					out<=243;
				end
				if(in == 1) begin
					state<=800;
					out<=244;
				end
				if(in == 2) begin
					state<=3697;
					out<=245;
				end
				if(in == 3) begin
					state<=5685;
					out<=246;
				end
				if(in == 4) begin
					state<=1796;
					out<=247;
				end
			end
			7576: begin
				if(in == 0) begin
					state<=7587;
					out<=248;
				end
				if(in == 1) begin
					state<=800;
					out<=249;
				end
				if(in == 2) begin
					state<=3698;
					out<=250;
				end
				if(in == 3) begin
					state<=5686;
					out<=251;
				end
				if(in == 4) begin
					state<=1797;
					out<=252;
				end
			end
			7577: begin
				if(in == 0) begin
					state<=7578;
					out<=253;
				end
				if(in == 1) begin
					state<=800;
					out<=254;
				end
				if(in == 2) begin
					state<=3689;
					out<=255;
				end
				if(in == 3) begin
					state<=5677;
					out<=0;
				end
				if(in == 4) begin
					state<=1788;
					out<=1;
				end
			end
			7578: begin
				if(in == 0) begin
					state<=7589;
					out<=2;
				end
				if(in == 1) begin
					state<=800;
					out<=3;
				end
				if(in == 2) begin
					state<=3700;
					out<=4;
				end
				if(in == 3) begin
					state<=5688;
					out<=5;
				end
				if(in == 4) begin
					state<=1799;
					out<=6;
				end
			end
			7579: begin
				if(in == 0) begin
					state<=7590;
					out<=7;
				end
				if(in == 1) begin
					state<=800;
					out<=8;
				end
				if(in == 2) begin
					state<=3701;
					out<=9;
				end
				if(in == 3) begin
					state<=5689;
					out<=10;
				end
				if(in == 4) begin
					state<=1800;
					out<=11;
				end
			end
			7580: begin
				if(in == 0) begin
					state<=7591;
					out<=12;
				end
				if(in == 1) begin
					state<=800;
					out<=13;
				end
				if(in == 2) begin
					state<=3702;
					out<=14;
				end
				if(in == 3) begin
					state<=5690;
					out<=15;
				end
				if(in == 4) begin
					state<=1801;
					out<=16;
				end
			end
			7581: begin
				if(in == 0) begin
					state<=7592;
					out<=17;
				end
				if(in == 1) begin
					state<=800;
					out<=18;
				end
				if(in == 2) begin
					state<=3703;
					out<=19;
				end
				if(in == 3) begin
					state<=5691;
					out<=20;
				end
				if(in == 4) begin
					state<=1802;
					out<=21;
				end
			end
			7582: begin
				if(in == 0) begin
					state<=7593;
					out<=22;
				end
				if(in == 1) begin
					state<=800;
					out<=23;
				end
				if(in == 2) begin
					state<=3704;
					out<=24;
				end
				if(in == 3) begin
					state<=5692;
					out<=25;
				end
				if(in == 4) begin
					state<=1803;
					out<=26;
				end
			end
			7583: begin
				if(in == 0) begin
					state<=7594;
					out<=27;
				end
				if(in == 1) begin
					state<=800;
					out<=28;
				end
				if(in == 2) begin
					state<=3705;
					out<=29;
				end
				if(in == 3) begin
					state<=5693;
					out<=30;
				end
				if(in == 4) begin
					state<=1804;
					out<=31;
				end
			end
			7584: begin
				if(in == 0) begin
					state<=7595;
					out<=32;
				end
				if(in == 1) begin
					state<=800;
					out<=33;
				end
				if(in == 2) begin
					state<=3706;
					out<=34;
				end
				if(in == 3) begin
					state<=5694;
					out<=35;
				end
				if(in == 4) begin
					state<=1805;
					out<=36;
				end
			end
			7585: begin
				if(in == 0) begin
					state<=7596;
					out<=37;
				end
				if(in == 1) begin
					state<=800;
					out<=38;
				end
				if(in == 2) begin
					state<=3707;
					out<=39;
				end
				if(in == 3) begin
					state<=5695;
					out<=40;
				end
				if(in == 4) begin
					state<=1806;
					out<=41;
				end
			end
			7586: begin
				if(in == 0) begin
					state<=7597;
					out<=42;
				end
				if(in == 1) begin
					state<=800;
					out<=43;
				end
				if(in == 2) begin
					state<=3708;
					out<=44;
				end
				if(in == 3) begin
					state<=5696;
					out<=45;
				end
				if(in == 4) begin
					state<=1807;
					out<=46;
				end
			end
			7587: begin
				if(in == 0) begin
					state<=7588;
					out<=47;
				end
				if(in == 1) begin
					state<=800;
					out<=48;
				end
				if(in == 2) begin
					state<=3699;
					out<=49;
				end
				if(in == 3) begin
					state<=5687;
					out<=50;
				end
				if(in == 4) begin
					state<=1798;
					out<=51;
				end
			end
			7588: begin
				if(in == 0) begin
					state<=7599;
					out<=52;
				end
				if(in == 1) begin
					state<=800;
					out<=53;
				end
				if(in == 2) begin
					state<=3710;
					out<=54;
				end
				if(in == 3) begin
					state<=5698;
					out<=55;
				end
				if(in == 4) begin
					state<=1809;
					out<=56;
				end
			end
			7589: begin
				if(in == 0) begin
					state<=7600;
					out<=57;
				end
				if(in == 1) begin
					state<=800;
					out<=58;
				end
				if(in == 2) begin
					state<=3711;
					out<=59;
				end
				if(in == 3) begin
					state<=5699;
					out<=60;
				end
				if(in == 4) begin
					state<=1810;
					out<=61;
				end
			end
			7590: begin
				if(in == 0) begin
					state<=7601;
					out<=62;
				end
				if(in == 1) begin
					state<=800;
					out<=63;
				end
				if(in == 2) begin
					state<=3712;
					out<=64;
				end
				if(in == 3) begin
					state<=5700;
					out<=65;
				end
				if(in == 4) begin
					state<=1811;
					out<=66;
				end
			end
			7591: begin
				if(in == 0) begin
					state<=7602;
					out<=67;
				end
				if(in == 1) begin
					state<=800;
					out<=68;
				end
				if(in == 2) begin
					state<=3713;
					out<=69;
				end
				if(in == 3) begin
					state<=5701;
					out<=70;
				end
				if(in == 4) begin
					state<=1812;
					out<=71;
				end
			end
			7592: begin
				if(in == 0) begin
					state<=7603;
					out<=72;
				end
				if(in == 1) begin
					state<=800;
					out<=73;
				end
				if(in == 2) begin
					state<=3714;
					out<=74;
				end
				if(in == 3) begin
					state<=5702;
					out<=75;
				end
				if(in == 4) begin
					state<=1813;
					out<=76;
				end
			end
			7593: begin
				if(in == 0) begin
					state<=7604;
					out<=77;
				end
				if(in == 1) begin
					state<=800;
					out<=78;
				end
				if(in == 2) begin
					state<=3715;
					out<=79;
				end
				if(in == 3) begin
					state<=5703;
					out<=80;
				end
				if(in == 4) begin
					state<=1814;
					out<=81;
				end
			end
			7594: begin
				if(in == 0) begin
					state<=7605;
					out<=82;
				end
				if(in == 1) begin
					state<=800;
					out<=83;
				end
				if(in == 2) begin
					state<=3716;
					out<=84;
				end
				if(in == 3) begin
					state<=5704;
					out<=85;
				end
				if(in == 4) begin
					state<=1815;
					out<=86;
				end
			end
			7595: begin
				if(in == 0) begin
					state<=7606;
					out<=87;
				end
				if(in == 1) begin
					state<=800;
					out<=88;
				end
				if(in == 2) begin
					state<=3717;
					out<=89;
				end
				if(in == 3) begin
					state<=5705;
					out<=90;
				end
				if(in == 4) begin
					state<=1816;
					out<=91;
				end
			end
			7596: begin
				if(in == 0) begin
					state<=7607;
					out<=92;
				end
				if(in == 1) begin
					state<=800;
					out<=93;
				end
				if(in == 2) begin
					state<=3718;
					out<=94;
				end
				if(in == 3) begin
					state<=5706;
					out<=95;
				end
				if(in == 4) begin
					state<=1817;
					out<=96;
				end
			end
			7597: begin
				if(in == 0) begin
					state<=7598;
					out<=97;
				end
				if(in == 1) begin
					state<=800;
					out<=98;
				end
				if(in == 2) begin
					state<=3709;
					out<=99;
				end
				if(in == 3) begin
					state<=5697;
					out<=100;
				end
				if(in == 4) begin
					state<=1808;
					out<=101;
				end
			end
			7598: begin
				if(in == 0) begin
					state<=7609;
					out<=102;
				end
				if(in == 1) begin
					state<=800;
					out<=103;
				end
				if(in == 2) begin
					state<=3720;
					out<=104;
				end
				if(in == 3) begin
					state<=5708;
					out<=105;
				end
				if(in == 4) begin
					state<=1819;
					out<=106;
				end
			end
			7599: begin
				if(in == 0) begin
					state<=7610;
					out<=107;
				end
				if(in == 1) begin
					state<=800;
					out<=108;
				end
				if(in == 2) begin
					state<=3721;
					out<=109;
				end
				if(in == 3) begin
					state<=5709;
					out<=110;
				end
				if(in == 4) begin
					state<=1820;
					out<=111;
				end
			end
			7600: begin
				if(in == 0) begin
					state<=7611;
					out<=112;
				end
				if(in == 1) begin
					state<=800;
					out<=113;
				end
				if(in == 2) begin
					state<=3722;
					out<=114;
				end
				if(in == 3) begin
					state<=5710;
					out<=115;
				end
				if(in == 4) begin
					state<=1821;
					out<=116;
				end
			end
			7601: begin
				if(in == 0) begin
					state<=7612;
					out<=117;
				end
				if(in == 1) begin
					state<=800;
					out<=118;
				end
				if(in == 2) begin
					state<=3723;
					out<=119;
				end
				if(in == 3) begin
					state<=5711;
					out<=120;
				end
				if(in == 4) begin
					state<=1822;
					out<=121;
				end
			end
			7602: begin
				if(in == 0) begin
					state<=7613;
					out<=122;
				end
				if(in == 1) begin
					state<=800;
					out<=123;
				end
				if(in == 2) begin
					state<=3724;
					out<=124;
				end
				if(in == 3) begin
					state<=5712;
					out<=125;
				end
				if(in == 4) begin
					state<=1823;
					out<=126;
				end
			end
			7603: begin
				if(in == 0) begin
					state<=7614;
					out<=127;
				end
				if(in == 1) begin
					state<=800;
					out<=128;
				end
				if(in == 2) begin
					state<=3725;
					out<=129;
				end
				if(in == 3) begin
					state<=5713;
					out<=130;
				end
				if(in == 4) begin
					state<=1824;
					out<=131;
				end
			end
			7604: begin
				if(in == 0) begin
					state<=7615;
					out<=132;
				end
				if(in == 1) begin
					state<=800;
					out<=133;
				end
				if(in == 2) begin
					state<=3726;
					out<=134;
				end
				if(in == 3) begin
					state<=5714;
					out<=135;
				end
				if(in == 4) begin
					state<=1825;
					out<=136;
				end
			end
			7605: begin
				if(in == 0) begin
					state<=7616;
					out<=137;
				end
				if(in == 1) begin
					state<=800;
					out<=138;
				end
				if(in == 2) begin
					state<=3727;
					out<=139;
				end
				if(in == 3) begin
					state<=5715;
					out<=140;
				end
				if(in == 4) begin
					state<=1826;
					out<=141;
				end
			end
			7606: begin
				if(in == 0) begin
					state<=7617;
					out<=142;
				end
				if(in == 1) begin
					state<=800;
					out<=143;
				end
				if(in == 2) begin
					state<=3728;
					out<=144;
				end
				if(in == 3) begin
					state<=5716;
					out<=145;
				end
				if(in == 4) begin
					state<=1827;
					out<=146;
				end
			end
			7607: begin
				if(in == 0) begin
					state<=7608;
					out<=147;
				end
				if(in == 1) begin
					state<=800;
					out<=148;
				end
				if(in == 2) begin
					state<=3719;
					out<=149;
				end
				if(in == 3) begin
					state<=5707;
					out<=150;
				end
				if(in == 4) begin
					state<=1818;
					out<=151;
				end
			end
			7608: begin
				if(in == 0) begin
					state<=7619;
					out<=152;
				end
				if(in == 1) begin
					state<=800;
					out<=153;
				end
				if(in == 2) begin
					state<=3730;
					out<=154;
				end
				if(in == 3) begin
					state<=5718;
					out<=155;
				end
				if(in == 4) begin
					state<=1829;
					out<=156;
				end
			end
			7609: begin
				if(in == 0) begin
					state<=7620;
					out<=157;
				end
				if(in == 1) begin
					state<=800;
					out<=158;
				end
				if(in == 2) begin
					state<=3731;
					out<=159;
				end
				if(in == 3) begin
					state<=5719;
					out<=160;
				end
				if(in == 4) begin
					state<=1830;
					out<=161;
				end
			end
			7610: begin
				if(in == 0) begin
					state<=7621;
					out<=162;
				end
				if(in == 1) begin
					state<=800;
					out<=163;
				end
				if(in == 2) begin
					state<=3732;
					out<=164;
				end
				if(in == 3) begin
					state<=5720;
					out<=165;
				end
				if(in == 4) begin
					state<=1831;
					out<=166;
				end
			end
			7611: begin
				if(in == 0) begin
					state<=7622;
					out<=167;
				end
				if(in == 1) begin
					state<=800;
					out<=168;
				end
				if(in == 2) begin
					state<=3733;
					out<=169;
				end
				if(in == 3) begin
					state<=5721;
					out<=170;
				end
				if(in == 4) begin
					state<=1832;
					out<=171;
				end
			end
			7612: begin
				if(in == 0) begin
					state<=7623;
					out<=172;
				end
				if(in == 1) begin
					state<=800;
					out<=173;
				end
				if(in == 2) begin
					state<=3734;
					out<=174;
				end
				if(in == 3) begin
					state<=5722;
					out<=175;
				end
				if(in == 4) begin
					state<=1833;
					out<=176;
				end
			end
			7613: begin
				if(in == 0) begin
					state<=7624;
					out<=177;
				end
				if(in == 1) begin
					state<=800;
					out<=178;
				end
				if(in == 2) begin
					state<=3735;
					out<=179;
				end
				if(in == 3) begin
					state<=5723;
					out<=180;
				end
				if(in == 4) begin
					state<=1834;
					out<=181;
				end
			end
			7614: begin
				if(in == 0) begin
					state<=7625;
					out<=182;
				end
				if(in == 1) begin
					state<=800;
					out<=183;
				end
				if(in == 2) begin
					state<=3736;
					out<=184;
				end
				if(in == 3) begin
					state<=5724;
					out<=185;
				end
				if(in == 4) begin
					state<=1835;
					out<=186;
				end
			end
			7615: begin
				if(in == 0) begin
					state<=7626;
					out<=187;
				end
				if(in == 1) begin
					state<=800;
					out<=188;
				end
				if(in == 2) begin
					state<=3737;
					out<=189;
				end
				if(in == 3) begin
					state<=5725;
					out<=190;
				end
				if(in == 4) begin
					state<=1836;
					out<=191;
				end
			end
			7616: begin
				if(in == 0) begin
					state<=7627;
					out<=192;
				end
				if(in == 1) begin
					state<=800;
					out<=193;
				end
				if(in == 2) begin
					state<=3738;
					out<=194;
				end
				if(in == 3) begin
					state<=5726;
					out<=195;
				end
				if(in == 4) begin
					state<=1837;
					out<=196;
				end
			end
			7617: begin
				if(in == 0) begin
					state<=7618;
					out<=197;
				end
				if(in == 1) begin
					state<=800;
					out<=198;
				end
				if(in == 2) begin
					state<=3729;
					out<=199;
				end
				if(in == 3) begin
					state<=5717;
					out<=200;
				end
				if(in == 4) begin
					state<=1828;
					out<=201;
				end
			end
			7618: begin
				if(in == 0) begin
					state<=7629;
					out<=202;
				end
				if(in == 1) begin
					state<=800;
					out<=203;
				end
				if(in == 2) begin
					state<=3740;
					out<=204;
				end
				if(in == 3) begin
					state<=5728;
					out<=205;
				end
				if(in == 4) begin
					state<=1839;
					out<=206;
				end
			end
			7619: begin
				if(in == 0) begin
					state<=7630;
					out<=207;
				end
				if(in == 1) begin
					state<=800;
					out<=208;
				end
				if(in == 2) begin
					state<=3741;
					out<=209;
				end
				if(in == 3) begin
					state<=5729;
					out<=210;
				end
				if(in == 4) begin
					state<=1840;
					out<=211;
				end
			end
			7620: begin
				if(in == 0) begin
					state<=7631;
					out<=212;
				end
				if(in == 1) begin
					state<=800;
					out<=213;
				end
				if(in == 2) begin
					state<=3742;
					out<=214;
				end
				if(in == 3) begin
					state<=5730;
					out<=215;
				end
				if(in == 4) begin
					state<=1841;
					out<=216;
				end
			end
			7621: begin
				if(in == 0) begin
					state<=7632;
					out<=217;
				end
				if(in == 1) begin
					state<=800;
					out<=218;
				end
				if(in == 2) begin
					state<=3743;
					out<=219;
				end
				if(in == 3) begin
					state<=5731;
					out<=220;
				end
				if(in == 4) begin
					state<=1842;
					out<=221;
				end
			end
			7622: begin
				if(in == 0) begin
					state<=7633;
					out<=222;
				end
				if(in == 1) begin
					state<=800;
					out<=223;
				end
				if(in == 2) begin
					state<=3744;
					out<=224;
				end
				if(in == 3) begin
					state<=5732;
					out<=225;
				end
				if(in == 4) begin
					state<=1843;
					out<=226;
				end
			end
			7623: begin
				if(in == 0) begin
					state<=7634;
					out<=227;
				end
				if(in == 1) begin
					state<=800;
					out<=228;
				end
				if(in == 2) begin
					state<=3745;
					out<=229;
				end
				if(in == 3) begin
					state<=5733;
					out<=230;
				end
				if(in == 4) begin
					state<=1844;
					out<=231;
				end
			end
			7624: begin
				if(in == 0) begin
					state<=7635;
					out<=232;
				end
				if(in == 1) begin
					state<=800;
					out<=233;
				end
				if(in == 2) begin
					state<=3746;
					out<=234;
				end
				if(in == 3) begin
					state<=5734;
					out<=235;
				end
				if(in == 4) begin
					state<=1845;
					out<=236;
				end
			end
			7625: begin
				if(in == 0) begin
					state<=7636;
					out<=237;
				end
				if(in == 1) begin
					state<=800;
					out<=238;
				end
				if(in == 2) begin
					state<=3747;
					out<=239;
				end
				if(in == 3) begin
					state<=5735;
					out<=240;
				end
				if(in == 4) begin
					state<=1846;
					out<=241;
				end
			end
			7626: begin
				if(in == 0) begin
					state<=7637;
					out<=242;
				end
				if(in == 1) begin
					state<=800;
					out<=243;
				end
				if(in == 2) begin
					state<=3748;
					out<=244;
				end
				if(in == 3) begin
					state<=5736;
					out<=245;
				end
				if(in == 4) begin
					state<=1847;
					out<=246;
				end
			end
			7627: begin
				if(in == 0) begin
					state<=7628;
					out<=247;
				end
				if(in == 1) begin
					state<=800;
					out<=248;
				end
				if(in == 2) begin
					state<=3739;
					out<=249;
				end
				if(in == 3) begin
					state<=5727;
					out<=250;
				end
				if(in == 4) begin
					state<=1838;
					out<=251;
				end
			end
			7628: begin
				if(in == 0) begin
					state<=7639;
					out<=252;
				end
				if(in == 1) begin
					state<=800;
					out<=253;
				end
				if(in == 2) begin
					state<=3750;
					out<=254;
				end
				if(in == 3) begin
					state<=5738;
					out<=255;
				end
				if(in == 4) begin
					state<=1849;
					out<=0;
				end
			end
			7629: begin
				if(in == 0) begin
					state<=7640;
					out<=1;
				end
				if(in == 1) begin
					state<=800;
					out<=2;
				end
				if(in == 2) begin
					state<=3751;
					out<=3;
				end
				if(in == 3) begin
					state<=5739;
					out<=4;
				end
				if(in == 4) begin
					state<=1850;
					out<=5;
				end
			end
			7630: begin
				if(in == 0) begin
					state<=7641;
					out<=6;
				end
				if(in == 1) begin
					state<=800;
					out<=7;
				end
				if(in == 2) begin
					state<=3752;
					out<=8;
				end
				if(in == 3) begin
					state<=5740;
					out<=9;
				end
				if(in == 4) begin
					state<=1851;
					out<=10;
				end
			end
			7631: begin
				if(in == 0) begin
					state<=7642;
					out<=11;
				end
				if(in == 1) begin
					state<=800;
					out<=12;
				end
				if(in == 2) begin
					state<=3753;
					out<=13;
				end
				if(in == 3) begin
					state<=5741;
					out<=14;
				end
				if(in == 4) begin
					state<=1852;
					out<=15;
				end
			end
			7632: begin
				if(in == 0) begin
					state<=7643;
					out<=16;
				end
				if(in == 1) begin
					state<=800;
					out<=17;
				end
				if(in == 2) begin
					state<=3754;
					out<=18;
				end
				if(in == 3) begin
					state<=5742;
					out<=19;
				end
				if(in == 4) begin
					state<=1853;
					out<=20;
				end
			end
			7633: begin
				if(in == 0) begin
					state<=7644;
					out<=21;
				end
				if(in == 1) begin
					state<=800;
					out<=22;
				end
				if(in == 2) begin
					state<=3755;
					out<=23;
				end
				if(in == 3) begin
					state<=5743;
					out<=24;
				end
				if(in == 4) begin
					state<=1854;
					out<=25;
				end
			end
			7634: begin
				if(in == 0) begin
					state<=7645;
					out<=26;
				end
				if(in == 1) begin
					state<=800;
					out<=27;
				end
				if(in == 2) begin
					state<=3756;
					out<=28;
				end
				if(in == 3) begin
					state<=5744;
					out<=29;
				end
				if(in == 4) begin
					state<=1855;
					out<=30;
				end
			end
			7635: begin
				if(in == 0) begin
					state<=7646;
					out<=31;
				end
				if(in == 1) begin
					state<=800;
					out<=32;
				end
				if(in == 2) begin
					state<=3757;
					out<=33;
				end
				if(in == 3) begin
					state<=5745;
					out<=34;
				end
				if(in == 4) begin
					state<=1856;
					out<=35;
				end
			end
			7636: begin
				if(in == 0) begin
					state<=7647;
					out<=36;
				end
				if(in == 1) begin
					state<=800;
					out<=37;
				end
				if(in == 2) begin
					state<=3758;
					out<=38;
				end
				if(in == 3) begin
					state<=5746;
					out<=39;
				end
				if(in == 4) begin
					state<=1857;
					out<=40;
				end
			end
			7637: begin
				if(in == 0) begin
					state<=7638;
					out<=41;
				end
				if(in == 1) begin
					state<=800;
					out<=42;
				end
				if(in == 2) begin
					state<=3749;
					out<=43;
				end
				if(in == 3) begin
					state<=5737;
					out<=44;
				end
				if(in == 4) begin
					state<=1848;
					out<=45;
				end
			end
			7638: begin
				if(in == 0) begin
					state<=7649;
					out<=46;
				end
				if(in == 1) begin
					state<=800;
					out<=47;
				end
				if(in == 2) begin
					state<=3760;
					out<=48;
				end
				if(in == 3) begin
					state<=5748;
					out<=49;
				end
				if(in == 4) begin
					state<=1859;
					out<=50;
				end
			end
			7639: begin
				if(in == 0) begin
					state<=7650;
					out<=51;
				end
				if(in == 1) begin
					state<=800;
					out<=52;
				end
				if(in == 2) begin
					state<=3761;
					out<=53;
				end
				if(in == 3) begin
					state<=5749;
					out<=54;
				end
				if(in == 4) begin
					state<=1860;
					out<=55;
				end
			end
			7640: begin
				if(in == 0) begin
					state<=7651;
					out<=56;
				end
				if(in == 1) begin
					state<=800;
					out<=57;
				end
				if(in == 2) begin
					state<=3762;
					out<=58;
				end
				if(in == 3) begin
					state<=5750;
					out<=59;
				end
				if(in == 4) begin
					state<=1861;
					out<=60;
				end
			end
			7641: begin
				if(in == 0) begin
					state<=7652;
					out<=61;
				end
				if(in == 1) begin
					state<=800;
					out<=62;
				end
				if(in == 2) begin
					state<=3763;
					out<=63;
				end
				if(in == 3) begin
					state<=5751;
					out<=64;
				end
				if(in == 4) begin
					state<=1862;
					out<=65;
				end
			end
			7642: begin
				if(in == 0) begin
					state<=7653;
					out<=66;
				end
				if(in == 1) begin
					state<=800;
					out<=67;
				end
				if(in == 2) begin
					state<=3764;
					out<=68;
				end
				if(in == 3) begin
					state<=5752;
					out<=69;
				end
				if(in == 4) begin
					state<=1863;
					out<=70;
				end
			end
			7643: begin
				if(in == 0) begin
					state<=7654;
					out<=71;
				end
				if(in == 1) begin
					state<=800;
					out<=72;
				end
				if(in == 2) begin
					state<=3765;
					out<=73;
				end
				if(in == 3) begin
					state<=5753;
					out<=74;
				end
				if(in == 4) begin
					state<=1864;
					out<=75;
				end
			end
			7644: begin
				if(in == 0) begin
					state<=7655;
					out<=76;
				end
				if(in == 1) begin
					state<=800;
					out<=77;
				end
				if(in == 2) begin
					state<=3766;
					out<=78;
				end
				if(in == 3) begin
					state<=5754;
					out<=79;
				end
				if(in == 4) begin
					state<=1865;
					out<=80;
				end
			end
			7645: begin
				if(in == 0) begin
					state<=7656;
					out<=81;
				end
				if(in == 1) begin
					state<=800;
					out<=82;
				end
				if(in == 2) begin
					state<=3767;
					out<=83;
				end
				if(in == 3) begin
					state<=5755;
					out<=84;
				end
				if(in == 4) begin
					state<=1866;
					out<=85;
				end
			end
			7646: begin
				if(in == 0) begin
					state<=7657;
					out<=86;
				end
				if(in == 1) begin
					state<=800;
					out<=87;
				end
				if(in == 2) begin
					state<=3768;
					out<=88;
				end
				if(in == 3) begin
					state<=5756;
					out<=89;
				end
				if(in == 4) begin
					state<=1867;
					out<=90;
				end
			end
			7647: begin
				if(in == 0) begin
					state<=7648;
					out<=91;
				end
				if(in == 1) begin
					state<=800;
					out<=92;
				end
				if(in == 2) begin
					state<=3759;
					out<=93;
				end
				if(in == 3) begin
					state<=5747;
					out<=94;
				end
				if(in == 4) begin
					state<=1858;
					out<=95;
				end
			end
			7648: begin
				if(in == 0) begin
					state<=7659;
					out<=96;
				end
				if(in == 1) begin
					state<=800;
					out<=97;
				end
				if(in == 2) begin
					state<=3770;
					out<=98;
				end
				if(in == 3) begin
					state<=5758;
					out<=99;
				end
				if(in == 4) begin
					state<=1869;
					out<=100;
				end
			end
			7649: begin
				if(in == 0) begin
					state<=7660;
					out<=101;
				end
				if(in == 1) begin
					state<=800;
					out<=102;
				end
				if(in == 2) begin
					state<=3771;
					out<=103;
				end
				if(in == 3) begin
					state<=5759;
					out<=104;
				end
				if(in == 4) begin
					state<=1870;
					out<=105;
				end
			end
			7650: begin
				if(in == 0) begin
					state<=7661;
					out<=106;
				end
				if(in == 1) begin
					state<=800;
					out<=107;
				end
				if(in == 2) begin
					state<=3772;
					out<=108;
				end
				if(in == 3) begin
					state<=5760;
					out<=109;
				end
				if(in == 4) begin
					state<=1871;
					out<=110;
				end
			end
			7651: begin
				if(in == 0) begin
					state<=7662;
					out<=111;
				end
				if(in == 1) begin
					state<=800;
					out<=112;
				end
				if(in == 2) begin
					state<=3773;
					out<=113;
				end
				if(in == 3) begin
					state<=5761;
					out<=114;
				end
				if(in == 4) begin
					state<=1872;
					out<=115;
				end
			end
			7652: begin
				if(in == 0) begin
					state<=7663;
					out<=116;
				end
				if(in == 1) begin
					state<=800;
					out<=117;
				end
				if(in == 2) begin
					state<=3774;
					out<=118;
				end
				if(in == 3) begin
					state<=5762;
					out<=119;
				end
				if(in == 4) begin
					state<=1873;
					out<=120;
				end
			end
			7653: begin
				if(in == 0) begin
					state<=7664;
					out<=121;
				end
				if(in == 1) begin
					state<=800;
					out<=122;
				end
				if(in == 2) begin
					state<=3775;
					out<=123;
				end
				if(in == 3) begin
					state<=5763;
					out<=124;
				end
				if(in == 4) begin
					state<=1874;
					out<=125;
				end
			end
			7654: begin
				if(in == 0) begin
					state<=7665;
					out<=126;
				end
				if(in == 1) begin
					state<=800;
					out<=127;
				end
				if(in == 2) begin
					state<=3776;
					out<=128;
				end
				if(in == 3) begin
					state<=5764;
					out<=129;
				end
				if(in == 4) begin
					state<=1875;
					out<=130;
				end
			end
			7655: begin
				if(in == 0) begin
					state<=7666;
					out<=131;
				end
				if(in == 1) begin
					state<=800;
					out<=132;
				end
				if(in == 2) begin
					state<=3777;
					out<=133;
				end
				if(in == 3) begin
					state<=5765;
					out<=134;
				end
				if(in == 4) begin
					state<=1876;
					out<=135;
				end
			end
			7656: begin
				if(in == 0) begin
					state<=7667;
					out<=136;
				end
				if(in == 1) begin
					state<=800;
					out<=137;
				end
				if(in == 2) begin
					state<=3778;
					out<=138;
				end
				if(in == 3) begin
					state<=5766;
					out<=139;
				end
				if(in == 4) begin
					state<=1877;
					out<=140;
				end
			end
			7657: begin
				if(in == 0) begin
					state<=7658;
					out<=141;
				end
				if(in == 1) begin
					state<=800;
					out<=142;
				end
				if(in == 2) begin
					state<=3769;
					out<=143;
				end
				if(in == 3) begin
					state<=5757;
					out<=144;
				end
				if(in == 4) begin
					state<=1868;
					out<=145;
				end
			end
			7658: begin
				if(in == 0) begin
					state<=7669;
					out<=146;
				end
				if(in == 1) begin
					state<=800;
					out<=147;
				end
				if(in == 2) begin
					state<=3780;
					out<=148;
				end
				if(in == 3) begin
					state<=5768;
					out<=149;
				end
				if(in == 4) begin
					state<=1879;
					out<=150;
				end
			end
			7659: begin
				if(in == 0) begin
					state<=7670;
					out<=151;
				end
				if(in == 1) begin
					state<=800;
					out<=152;
				end
				if(in == 2) begin
					state<=3781;
					out<=153;
				end
				if(in == 3) begin
					state<=5769;
					out<=154;
				end
				if(in == 4) begin
					state<=1880;
					out<=155;
				end
			end
			7660: begin
				if(in == 0) begin
					state<=7671;
					out<=156;
				end
				if(in == 1) begin
					state<=800;
					out<=157;
				end
				if(in == 2) begin
					state<=3782;
					out<=158;
				end
				if(in == 3) begin
					state<=5770;
					out<=159;
				end
				if(in == 4) begin
					state<=1881;
					out<=160;
				end
			end
			7661: begin
				if(in == 0) begin
					state<=7672;
					out<=161;
				end
				if(in == 1) begin
					state<=800;
					out<=162;
				end
				if(in == 2) begin
					state<=3783;
					out<=163;
				end
				if(in == 3) begin
					state<=5771;
					out<=164;
				end
				if(in == 4) begin
					state<=1882;
					out<=165;
				end
			end
			7662: begin
				if(in == 0) begin
					state<=7673;
					out<=166;
				end
				if(in == 1) begin
					state<=800;
					out<=167;
				end
				if(in == 2) begin
					state<=3784;
					out<=168;
				end
				if(in == 3) begin
					state<=5772;
					out<=169;
				end
				if(in == 4) begin
					state<=1883;
					out<=170;
				end
			end
			7663: begin
				if(in == 0) begin
					state<=7674;
					out<=171;
				end
				if(in == 1) begin
					state<=800;
					out<=172;
				end
				if(in == 2) begin
					state<=3785;
					out<=173;
				end
				if(in == 3) begin
					state<=5773;
					out<=174;
				end
				if(in == 4) begin
					state<=1884;
					out<=175;
				end
			end
			7664: begin
				if(in == 0) begin
					state<=7675;
					out<=176;
				end
				if(in == 1) begin
					state<=800;
					out<=177;
				end
				if(in == 2) begin
					state<=3786;
					out<=178;
				end
				if(in == 3) begin
					state<=5774;
					out<=179;
				end
				if(in == 4) begin
					state<=1885;
					out<=180;
				end
			end
			7665: begin
				if(in == 0) begin
					state<=7676;
					out<=181;
				end
				if(in == 1) begin
					state<=800;
					out<=182;
				end
				if(in == 2) begin
					state<=3787;
					out<=183;
				end
				if(in == 3) begin
					state<=5775;
					out<=184;
				end
				if(in == 4) begin
					state<=1886;
					out<=185;
				end
			end
			7666: begin
				if(in == 0) begin
					state<=7677;
					out<=186;
				end
				if(in == 1) begin
					state<=800;
					out<=187;
				end
				if(in == 2) begin
					state<=3788;
					out<=188;
				end
				if(in == 3) begin
					state<=5776;
					out<=189;
				end
				if(in == 4) begin
					state<=1887;
					out<=190;
				end
			end
			7667: begin
				if(in == 0) begin
					state<=7668;
					out<=191;
				end
				if(in == 1) begin
					state<=800;
					out<=192;
				end
				if(in == 2) begin
					state<=3779;
					out<=193;
				end
				if(in == 3) begin
					state<=5767;
					out<=194;
				end
				if(in == 4) begin
					state<=1878;
					out<=195;
				end
			end
			7668: begin
				if(in == 0) begin
					state<=7679;
					out<=196;
				end
				if(in == 1) begin
					state<=800;
					out<=197;
				end
				if(in == 2) begin
					state<=3790;
					out<=198;
				end
				if(in == 3) begin
					state<=5778;
					out<=199;
				end
				if(in == 4) begin
					state<=1889;
					out<=200;
				end
			end
			7669: begin
				if(in == 0) begin
					state<=7680;
					out<=201;
				end
				if(in == 1) begin
					state<=800;
					out<=202;
				end
				if(in == 2) begin
					state<=3791;
					out<=203;
				end
				if(in == 3) begin
					state<=5779;
					out<=204;
				end
				if(in == 4) begin
					state<=1890;
					out<=205;
				end
			end
			7670: begin
				if(in == 0) begin
					state<=7681;
					out<=206;
				end
				if(in == 1) begin
					state<=800;
					out<=207;
				end
				if(in == 2) begin
					state<=3792;
					out<=208;
				end
				if(in == 3) begin
					state<=5780;
					out<=209;
				end
				if(in == 4) begin
					state<=1891;
					out<=210;
				end
			end
			7671: begin
				if(in == 0) begin
					state<=7682;
					out<=211;
				end
				if(in == 1) begin
					state<=800;
					out<=212;
				end
				if(in == 2) begin
					state<=3793;
					out<=213;
				end
				if(in == 3) begin
					state<=5781;
					out<=214;
				end
				if(in == 4) begin
					state<=1892;
					out<=215;
				end
			end
			7672: begin
				if(in == 0) begin
					state<=7683;
					out<=216;
				end
				if(in == 1) begin
					state<=800;
					out<=217;
				end
				if(in == 2) begin
					state<=3794;
					out<=218;
				end
				if(in == 3) begin
					state<=5782;
					out<=219;
				end
				if(in == 4) begin
					state<=1893;
					out<=220;
				end
			end
			7673: begin
				if(in == 0) begin
					state<=7684;
					out<=221;
				end
				if(in == 1) begin
					state<=800;
					out<=222;
				end
				if(in == 2) begin
					state<=3795;
					out<=223;
				end
				if(in == 3) begin
					state<=5783;
					out<=224;
				end
				if(in == 4) begin
					state<=1894;
					out<=225;
				end
			end
			7674: begin
				if(in == 0) begin
					state<=7685;
					out<=226;
				end
				if(in == 1) begin
					state<=800;
					out<=227;
				end
				if(in == 2) begin
					state<=3796;
					out<=228;
				end
				if(in == 3) begin
					state<=5784;
					out<=229;
				end
				if(in == 4) begin
					state<=1895;
					out<=230;
				end
			end
			7675: begin
				if(in == 0) begin
					state<=7686;
					out<=231;
				end
				if(in == 1) begin
					state<=800;
					out<=232;
				end
				if(in == 2) begin
					state<=3797;
					out<=233;
				end
				if(in == 3) begin
					state<=5785;
					out<=234;
				end
				if(in == 4) begin
					state<=1896;
					out<=235;
				end
			end
			7676: begin
				if(in == 0) begin
					state<=7687;
					out<=236;
				end
				if(in == 1) begin
					state<=800;
					out<=237;
				end
				if(in == 2) begin
					state<=3798;
					out<=238;
				end
				if(in == 3) begin
					state<=5786;
					out<=239;
				end
				if(in == 4) begin
					state<=1897;
					out<=240;
				end
			end
			7677: begin
				if(in == 0) begin
					state<=7678;
					out<=241;
				end
				if(in == 1) begin
					state<=800;
					out<=242;
				end
				if(in == 2) begin
					state<=3789;
					out<=243;
				end
				if(in == 3) begin
					state<=5777;
					out<=244;
				end
				if(in == 4) begin
					state<=1888;
					out<=245;
				end
			end
			7678: begin
				if(in == 0) begin
					state<=7689;
					out<=246;
				end
				if(in == 1) begin
					state<=800;
					out<=247;
				end
				if(in == 2) begin
					state<=3800;
					out<=248;
				end
				if(in == 3) begin
					state<=5788;
					out<=249;
				end
				if(in == 4) begin
					state<=1899;
					out<=250;
				end
			end
			7679: begin
				if(in == 0) begin
					state<=7690;
					out<=251;
				end
				if(in == 1) begin
					state<=800;
					out<=252;
				end
				if(in == 2) begin
					state<=3801;
					out<=253;
				end
				if(in == 3) begin
					state<=5789;
					out<=254;
				end
				if(in == 4) begin
					state<=1900;
					out<=255;
				end
			end
			7680: begin
				if(in == 0) begin
					state<=7691;
					out<=0;
				end
				if(in == 1) begin
					state<=800;
					out<=1;
				end
				if(in == 2) begin
					state<=3802;
					out<=2;
				end
				if(in == 3) begin
					state<=5790;
					out<=3;
				end
				if(in == 4) begin
					state<=1901;
					out<=4;
				end
			end
			7681: begin
				if(in == 0) begin
					state<=7692;
					out<=5;
				end
				if(in == 1) begin
					state<=800;
					out<=6;
				end
				if(in == 2) begin
					state<=3803;
					out<=7;
				end
				if(in == 3) begin
					state<=5791;
					out<=8;
				end
				if(in == 4) begin
					state<=1902;
					out<=9;
				end
			end
			7682: begin
				if(in == 0) begin
					state<=7693;
					out<=10;
				end
				if(in == 1) begin
					state<=800;
					out<=11;
				end
				if(in == 2) begin
					state<=3804;
					out<=12;
				end
				if(in == 3) begin
					state<=5792;
					out<=13;
				end
				if(in == 4) begin
					state<=1903;
					out<=14;
				end
			end
			7683: begin
				if(in == 0) begin
					state<=7694;
					out<=15;
				end
				if(in == 1) begin
					state<=800;
					out<=16;
				end
				if(in == 2) begin
					state<=3805;
					out<=17;
				end
				if(in == 3) begin
					state<=5793;
					out<=18;
				end
				if(in == 4) begin
					state<=1904;
					out<=19;
				end
			end
			7684: begin
				if(in == 0) begin
					state<=7695;
					out<=20;
				end
				if(in == 1) begin
					state<=800;
					out<=21;
				end
				if(in == 2) begin
					state<=3806;
					out<=22;
				end
				if(in == 3) begin
					state<=5794;
					out<=23;
				end
				if(in == 4) begin
					state<=1905;
					out<=24;
				end
			end
			7685: begin
				if(in == 0) begin
					state<=7696;
					out<=25;
				end
				if(in == 1) begin
					state<=800;
					out<=26;
				end
				if(in == 2) begin
					state<=3807;
					out<=27;
				end
				if(in == 3) begin
					state<=5795;
					out<=28;
				end
				if(in == 4) begin
					state<=1906;
					out<=29;
				end
			end
			7686: begin
				if(in == 0) begin
					state<=7697;
					out<=30;
				end
				if(in == 1) begin
					state<=800;
					out<=31;
				end
				if(in == 2) begin
					state<=3808;
					out<=32;
				end
				if(in == 3) begin
					state<=5796;
					out<=33;
				end
				if(in == 4) begin
					state<=1907;
					out<=34;
				end
			end
			7687: begin
				if(in == 0) begin
					state<=7688;
					out<=35;
				end
				if(in == 1) begin
					state<=800;
					out<=36;
				end
				if(in == 2) begin
					state<=3799;
					out<=37;
				end
				if(in == 3) begin
					state<=5787;
					out<=38;
				end
				if(in == 4) begin
					state<=1898;
					out<=39;
				end
			end
			7688: begin
				if(in == 0) begin
					state<=7699;
					out<=40;
				end
				if(in == 1) begin
					state<=800;
					out<=41;
				end
				if(in == 2) begin
					state<=3810;
					out<=42;
				end
				if(in == 3) begin
					state<=5798;
					out<=43;
				end
				if(in == 4) begin
					state<=1909;
					out<=44;
				end
			end
			7689: begin
				if(in == 0) begin
					state<=7700;
					out<=45;
				end
				if(in == 1) begin
					state<=800;
					out<=46;
				end
				if(in == 2) begin
					state<=3811;
					out<=47;
				end
				if(in == 3) begin
					state<=5799;
					out<=48;
				end
				if(in == 4) begin
					state<=1910;
					out<=49;
				end
			end
			7690: begin
				if(in == 0) begin
					state<=7701;
					out<=50;
				end
				if(in == 1) begin
					state<=800;
					out<=51;
				end
				if(in == 2) begin
					state<=3812;
					out<=52;
				end
				if(in == 3) begin
					state<=5800;
					out<=53;
				end
				if(in == 4) begin
					state<=1911;
					out<=54;
				end
			end
			7691: begin
				if(in == 0) begin
					state<=7702;
					out<=55;
				end
				if(in == 1) begin
					state<=800;
					out<=56;
				end
				if(in == 2) begin
					state<=3813;
					out<=57;
				end
				if(in == 3) begin
					state<=5801;
					out<=58;
				end
				if(in == 4) begin
					state<=1912;
					out<=59;
				end
			end
			7692: begin
				if(in == 0) begin
					state<=7703;
					out<=60;
				end
				if(in == 1) begin
					state<=800;
					out<=61;
				end
				if(in == 2) begin
					state<=3814;
					out<=62;
				end
				if(in == 3) begin
					state<=5802;
					out<=63;
				end
				if(in == 4) begin
					state<=1913;
					out<=64;
				end
			end
			7693: begin
				if(in == 0) begin
					state<=7704;
					out<=65;
				end
				if(in == 1) begin
					state<=800;
					out<=66;
				end
				if(in == 2) begin
					state<=3815;
					out<=67;
				end
				if(in == 3) begin
					state<=5803;
					out<=68;
				end
				if(in == 4) begin
					state<=1914;
					out<=69;
				end
			end
			7694: begin
				if(in == 0) begin
					state<=7705;
					out<=70;
				end
				if(in == 1) begin
					state<=800;
					out<=71;
				end
				if(in == 2) begin
					state<=3816;
					out<=72;
				end
				if(in == 3) begin
					state<=5804;
					out<=73;
				end
				if(in == 4) begin
					state<=1915;
					out<=74;
				end
			end
			7695: begin
				if(in == 0) begin
					state<=7706;
					out<=75;
				end
				if(in == 1) begin
					state<=800;
					out<=76;
				end
				if(in == 2) begin
					state<=3817;
					out<=77;
				end
				if(in == 3) begin
					state<=5805;
					out<=78;
				end
				if(in == 4) begin
					state<=1916;
					out<=79;
				end
			end
			7696: begin
				if(in == 0) begin
					state<=7707;
					out<=80;
				end
				if(in == 1) begin
					state<=800;
					out<=81;
				end
				if(in == 2) begin
					state<=3818;
					out<=82;
				end
				if(in == 3) begin
					state<=5806;
					out<=83;
				end
				if(in == 4) begin
					state<=1917;
					out<=84;
				end
			end
			7697: begin
				if(in == 0) begin
					state<=7698;
					out<=85;
				end
				if(in == 1) begin
					state<=800;
					out<=86;
				end
				if(in == 2) begin
					state<=3809;
					out<=87;
				end
				if(in == 3) begin
					state<=5797;
					out<=88;
				end
				if(in == 4) begin
					state<=1908;
					out<=89;
				end
			end
			7698: begin
				if(in == 0) begin
					state<=7709;
					out<=90;
				end
				if(in == 1) begin
					state<=800;
					out<=91;
				end
				if(in == 2) begin
					state<=3820;
					out<=92;
				end
				if(in == 3) begin
					state<=5808;
					out<=93;
				end
				if(in == 4) begin
					state<=1919;
					out<=94;
				end
			end
			7699: begin
				if(in == 0) begin
					state<=7710;
					out<=95;
				end
				if(in == 1) begin
					state<=800;
					out<=96;
				end
				if(in == 2) begin
					state<=3821;
					out<=97;
				end
				if(in == 3) begin
					state<=5809;
					out<=98;
				end
				if(in == 4) begin
					state<=1920;
					out<=99;
				end
			end
			7700: begin
				if(in == 0) begin
					state<=7711;
					out<=100;
				end
				if(in == 1) begin
					state<=800;
					out<=101;
				end
				if(in == 2) begin
					state<=3822;
					out<=102;
				end
				if(in == 3) begin
					state<=5810;
					out<=103;
				end
				if(in == 4) begin
					state<=1921;
					out<=104;
				end
			end
			7701: begin
				if(in == 0) begin
					state<=7712;
					out<=105;
				end
				if(in == 1) begin
					state<=800;
					out<=106;
				end
				if(in == 2) begin
					state<=3823;
					out<=107;
				end
				if(in == 3) begin
					state<=5811;
					out<=108;
				end
				if(in == 4) begin
					state<=1922;
					out<=109;
				end
			end
			7702: begin
				if(in == 0) begin
					state<=7713;
					out<=110;
				end
				if(in == 1) begin
					state<=800;
					out<=111;
				end
				if(in == 2) begin
					state<=3824;
					out<=112;
				end
				if(in == 3) begin
					state<=5812;
					out<=113;
				end
				if(in == 4) begin
					state<=1923;
					out<=114;
				end
			end
			7703: begin
				if(in == 0) begin
					state<=7714;
					out<=115;
				end
				if(in == 1) begin
					state<=800;
					out<=116;
				end
				if(in == 2) begin
					state<=3825;
					out<=117;
				end
				if(in == 3) begin
					state<=5813;
					out<=118;
				end
				if(in == 4) begin
					state<=1924;
					out<=119;
				end
			end
			7704: begin
				if(in == 0) begin
					state<=7715;
					out<=120;
				end
				if(in == 1) begin
					state<=800;
					out<=121;
				end
				if(in == 2) begin
					state<=3826;
					out<=122;
				end
				if(in == 3) begin
					state<=5814;
					out<=123;
				end
				if(in == 4) begin
					state<=1925;
					out<=124;
				end
			end
			7705: begin
				if(in == 0) begin
					state<=7716;
					out<=125;
				end
				if(in == 1) begin
					state<=800;
					out<=126;
				end
				if(in == 2) begin
					state<=3827;
					out<=127;
				end
				if(in == 3) begin
					state<=5815;
					out<=128;
				end
				if(in == 4) begin
					state<=1926;
					out<=129;
				end
			end
			7706: begin
				if(in == 0) begin
					state<=7717;
					out<=130;
				end
				if(in == 1) begin
					state<=800;
					out<=131;
				end
				if(in == 2) begin
					state<=3828;
					out<=132;
				end
				if(in == 3) begin
					state<=5816;
					out<=133;
				end
				if(in == 4) begin
					state<=1927;
					out<=134;
				end
			end
			7707: begin
				if(in == 0) begin
					state<=7708;
					out<=135;
				end
				if(in == 1) begin
					state<=800;
					out<=136;
				end
				if(in == 2) begin
					state<=3819;
					out<=137;
				end
				if(in == 3) begin
					state<=5807;
					out<=138;
				end
				if(in == 4) begin
					state<=1918;
					out<=139;
				end
			end
			7708: begin
				if(in == 0) begin
					state<=7719;
					out<=140;
				end
				if(in == 1) begin
					state<=800;
					out<=141;
				end
				if(in == 2) begin
					state<=3830;
					out<=142;
				end
				if(in == 3) begin
					state<=5818;
					out<=143;
				end
				if(in == 4) begin
					state<=1929;
					out<=144;
				end
			end
			7709: begin
				if(in == 0) begin
					state<=7720;
					out<=145;
				end
				if(in == 1) begin
					state<=800;
					out<=146;
				end
				if(in == 2) begin
					state<=3831;
					out<=147;
				end
				if(in == 3) begin
					state<=5819;
					out<=148;
				end
				if(in == 4) begin
					state<=1930;
					out<=149;
				end
			end
			7710: begin
				if(in == 0) begin
					state<=7721;
					out<=150;
				end
				if(in == 1) begin
					state<=800;
					out<=151;
				end
				if(in == 2) begin
					state<=3832;
					out<=152;
				end
				if(in == 3) begin
					state<=5820;
					out<=153;
				end
				if(in == 4) begin
					state<=1931;
					out<=154;
				end
			end
			7711: begin
				if(in == 0) begin
					state<=7722;
					out<=155;
				end
				if(in == 1) begin
					state<=800;
					out<=156;
				end
				if(in == 2) begin
					state<=3833;
					out<=157;
				end
				if(in == 3) begin
					state<=5821;
					out<=158;
				end
				if(in == 4) begin
					state<=1932;
					out<=159;
				end
			end
			7712: begin
				if(in == 0) begin
					state<=7723;
					out<=160;
				end
				if(in == 1) begin
					state<=800;
					out<=161;
				end
				if(in == 2) begin
					state<=3834;
					out<=162;
				end
				if(in == 3) begin
					state<=5822;
					out<=163;
				end
				if(in == 4) begin
					state<=1933;
					out<=164;
				end
			end
			7713: begin
				if(in == 0) begin
					state<=7724;
					out<=165;
				end
				if(in == 1) begin
					state<=800;
					out<=166;
				end
				if(in == 2) begin
					state<=3835;
					out<=167;
				end
				if(in == 3) begin
					state<=5823;
					out<=168;
				end
				if(in == 4) begin
					state<=1934;
					out<=169;
				end
			end
			7714: begin
				if(in == 0) begin
					state<=7725;
					out<=170;
				end
				if(in == 1) begin
					state<=800;
					out<=171;
				end
				if(in == 2) begin
					state<=3836;
					out<=172;
				end
				if(in == 3) begin
					state<=5824;
					out<=173;
				end
				if(in == 4) begin
					state<=1935;
					out<=174;
				end
			end
			7715: begin
				if(in == 0) begin
					state<=7726;
					out<=175;
				end
				if(in == 1) begin
					state<=800;
					out<=176;
				end
				if(in == 2) begin
					state<=3837;
					out<=177;
				end
				if(in == 3) begin
					state<=5825;
					out<=178;
				end
				if(in == 4) begin
					state<=1936;
					out<=179;
				end
			end
			7716: begin
				if(in == 0) begin
					state<=7727;
					out<=180;
				end
				if(in == 1) begin
					state<=800;
					out<=181;
				end
				if(in == 2) begin
					state<=3838;
					out<=182;
				end
				if(in == 3) begin
					state<=5826;
					out<=183;
				end
				if(in == 4) begin
					state<=1937;
					out<=184;
				end
			end
			7717: begin
				if(in == 0) begin
					state<=7718;
					out<=185;
				end
				if(in == 1) begin
					state<=800;
					out<=186;
				end
				if(in == 2) begin
					state<=3829;
					out<=187;
				end
				if(in == 3) begin
					state<=5817;
					out<=188;
				end
				if(in == 4) begin
					state<=1928;
					out<=189;
				end
			end
			7718: begin
				if(in == 0) begin
					state<=7729;
					out<=190;
				end
				if(in == 1) begin
					state<=800;
					out<=191;
				end
				if(in == 2) begin
					state<=3840;
					out<=192;
				end
				if(in == 3) begin
					state<=5828;
					out<=193;
				end
				if(in == 4) begin
					state<=1939;
					out<=194;
				end
			end
			7719: begin
				if(in == 0) begin
					state<=7730;
					out<=195;
				end
				if(in == 1) begin
					state<=800;
					out<=196;
				end
				if(in == 2) begin
					state<=3841;
					out<=197;
				end
				if(in == 3) begin
					state<=5829;
					out<=198;
				end
				if(in == 4) begin
					state<=1940;
					out<=199;
				end
			end
			7720: begin
				if(in == 0) begin
					state<=7731;
					out<=200;
				end
				if(in == 1) begin
					state<=800;
					out<=201;
				end
				if(in == 2) begin
					state<=3842;
					out<=202;
				end
				if(in == 3) begin
					state<=5830;
					out<=203;
				end
				if(in == 4) begin
					state<=1941;
					out<=204;
				end
			end
			7721: begin
				if(in == 0) begin
					state<=7732;
					out<=205;
				end
				if(in == 1) begin
					state<=800;
					out<=206;
				end
				if(in == 2) begin
					state<=3843;
					out<=207;
				end
				if(in == 3) begin
					state<=5831;
					out<=208;
				end
				if(in == 4) begin
					state<=1942;
					out<=209;
				end
			end
			7722: begin
				if(in == 0) begin
					state<=7733;
					out<=210;
				end
				if(in == 1) begin
					state<=800;
					out<=211;
				end
				if(in == 2) begin
					state<=3844;
					out<=212;
				end
				if(in == 3) begin
					state<=5832;
					out<=213;
				end
				if(in == 4) begin
					state<=1943;
					out<=214;
				end
			end
			7723: begin
				if(in == 0) begin
					state<=7734;
					out<=215;
				end
				if(in == 1) begin
					state<=800;
					out<=216;
				end
				if(in == 2) begin
					state<=3845;
					out<=217;
				end
				if(in == 3) begin
					state<=5833;
					out<=218;
				end
				if(in == 4) begin
					state<=1944;
					out<=219;
				end
			end
			7724: begin
				if(in == 0) begin
					state<=7735;
					out<=220;
				end
				if(in == 1) begin
					state<=800;
					out<=221;
				end
				if(in == 2) begin
					state<=3846;
					out<=222;
				end
				if(in == 3) begin
					state<=5834;
					out<=223;
				end
				if(in == 4) begin
					state<=1945;
					out<=224;
				end
			end
			7725: begin
				if(in == 0) begin
					state<=7736;
					out<=225;
				end
				if(in == 1) begin
					state<=800;
					out<=226;
				end
				if(in == 2) begin
					state<=3847;
					out<=227;
				end
				if(in == 3) begin
					state<=5835;
					out<=228;
				end
				if(in == 4) begin
					state<=1946;
					out<=229;
				end
			end
			7726: begin
				if(in == 0) begin
					state<=7737;
					out<=230;
				end
				if(in == 1) begin
					state<=800;
					out<=231;
				end
				if(in == 2) begin
					state<=3848;
					out<=232;
				end
				if(in == 3) begin
					state<=5836;
					out<=233;
				end
				if(in == 4) begin
					state<=1947;
					out<=234;
				end
			end
			7727: begin
				if(in == 0) begin
					state<=7728;
					out<=235;
				end
				if(in == 1) begin
					state<=800;
					out<=236;
				end
				if(in == 2) begin
					state<=3839;
					out<=237;
				end
				if(in == 3) begin
					state<=5827;
					out<=238;
				end
				if(in == 4) begin
					state<=1938;
					out<=239;
				end
			end
			7728: begin
				if(in == 0) begin
					state<=7739;
					out<=240;
				end
				if(in == 1) begin
					state<=800;
					out<=241;
				end
				if(in == 2) begin
					state<=3850;
					out<=242;
				end
				if(in == 3) begin
					state<=5838;
					out<=243;
				end
				if(in == 4) begin
					state<=1949;
					out<=244;
				end
			end
			7729: begin
				if(in == 0) begin
					state<=7740;
					out<=245;
				end
				if(in == 1) begin
					state<=800;
					out<=246;
				end
				if(in == 2) begin
					state<=3851;
					out<=247;
				end
				if(in == 3) begin
					state<=5839;
					out<=248;
				end
				if(in == 4) begin
					state<=1950;
					out<=249;
				end
			end
			7730: begin
				if(in == 0) begin
					state<=7741;
					out<=250;
				end
				if(in == 1) begin
					state<=800;
					out<=251;
				end
				if(in == 2) begin
					state<=3852;
					out<=252;
				end
				if(in == 3) begin
					state<=5840;
					out<=253;
				end
				if(in == 4) begin
					state<=1951;
					out<=254;
				end
			end
			7731: begin
				if(in == 0) begin
					state<=7742;
					out<=255;
				end
				if(in == 1) begin
					state<=800;
					out<=0;
				end
				if(in == 2) begin
					state<=3853;
					out<=1;
				end
				if(in == 3) begin
					state<=5841;
					out<=2;
				end
				if(in == 4) begin
					state<=1952;
					out<=3;
				end
			end
			7732: begin
				if(in == 0) begin
					state<=7743;
					out<=4;
				end
				if(in == 1) begin
					state<=800;
					out<=5;
				end
				if(in == 2) begin
					state<=3854;
					out<=6;
				end
				if(in == 3) begin
					state<=5842;
					out<=7;
				end
				if(in == 4) begin
					state<=1953;
					out<=8;
				end
			end
			7733: begin
				if(in == 0) begin
					state<=7744;
					out<=9;
				end
				if(in == 1) begin
					state<=800;
					out<=10;
				end
				if(in == 2) begin
					state<=3855;
					out<=11;
				end
				if(in == 3) begin
					state<=5843;
					out<=12;
				end
				if(in == 4) begin
					state<=1954;
					out<=13;
				end
			end
			7734: begin
				if(in == 0) begin
					state<=7745;
					out<=14;
				end
				if(in == 1) begin
					state<=800;
					out<=15;
				end
				if(in == 2) begin
					state<=3856;
					out<=16;
				end
				if(in == 3) begin
					state<=5844;
					out<=17;
				end
				if(in == 4) begin
					state<=1955;
					out<=18;
				end
			end
			7735: begin
				if(in == 0) begin
					state<=7746;
					out<=19;
				end
				if(in == 1) begin
					state<=800;
					out<=20;
				end
				if(in == 2) begin
					state<=3857;
					out<=21;
				end
				if(in == 3) begin
					state<=5845;
					out<=22;
				end
				if(in == 4) begin
					state<=1956;
					out<=23;
				end
			end
			7736: begin
				if(in == 0) begin
					state<=7747;
					out<=24;
				end
				if(in == 1) begin
					state<=800;
					out<=25;
				end
				if(in == 2) begin
					state<=3858;
					out<=26;
				end
				if(in == 3) begin
					state<=5846;
					out<=27;
				end
				if(in == 4) begin
					state<=1957;
					out<=28;
				end
			end
			7737: begin
				if(in == 0) begin
					state<=7738;
					out<=29;
				end
				if(in == 1) begin
					state<=800;
					out<=30;
				end
				if(in == 2) begin
					state<=3849;
					out<=31;
				end
				if(in == 3) begin
					state<=5837;
					out<=32;
				end
				if(in == 4) begin
					state<=1948;
					out<=33;
				end
			end
			7738: begin
				if(in == 0) begin
					state<=7749;
					out<=34;
				end
				if(in == 1) begin
					state<=800;
					out<=35;
				end
				if(in == 2) begin
					state<=3860;
					out<=36;
				end
				if(in == 3) begin
					state<=5848;
					out<=37;
				end
				if(in == 4) begin
					state<=1959;
					out<=38;
				end
			end
			7739: begin
				if(in == 0) begin
					state<=7750;
					out<=39;
				end
				if(in == 1) begin
					state<=800;
					out<=40;
				end
				if(in == 2) begin
					state<=3861;
					out<=41;
				end
				if(in == 3) begin
					state<=5849;
					out<=42;
				end
				if(in == 4) begin
					state<=1960;
					out<=43;
				end
			end
			7740: begin
				if(in == 0) begin
					state<=7751;
					out<=44;
				end
				if(in == 1) begin
					state<=800;
					out<=45;
				end
				if(in == 2) begin
					state<=3862;
					out<=46;
				end
				if(in == 3) begin
					state<=5850;
					out<=47;
				end
				if(in == 4) begin
					state<=1961;
					out<=48;
				end
			end
			7741: begin
				if(in == 0) begin
					state<=7752;
					out<=49;
				end
				if(in == 1) begin
					state<=800;
					out<=50;
				end
				if(in == 2) begin
					state<=3863;
					out<=51;
				end
				if(in == 3) begin
					state<=5851;
					out<=52;
				end
				if(in == 4) begin
					state<=1962;
					out<=53;
				end
			end
			7742: begin
				if(in == 0) begin
					state<=7753;
					out<=54;
				end
				if(in == 1) begin
					state<=800;
					out<=55;
				end
				if(in == 2) begin
					state<=3864;
					out<=56;
				end
				if(in == 3) begin
					state<=5852;
					out<=57;
				end
				if(in == 4) begin
					state<=1963;
					out<=58;
				end
			end
			7743: begin
				if(in == 0) begin
					state<=7754;
					out<=59;
				end
				if(in == 1) begin
					state<=800;
					out<=60;
				end
				if(in == 2) begin
					state<=3865;
					out<=61;
				end
				if(in == 3) begin
					state<=5853;
					out<=62;
				end
				if(in == 4) begin
					state<=1964;
					out<=63;
				end
			end
			7744: begin
				if(in == 0) begin
					state<=7755;
					out<=64;
				end
				if(in == 1) begin
					state<=800;
					out<=65;
				end
				if(in == 2) begin
					state<=3866;
					out<=66;
				end
				if(in == 3) begin
					state<=5854;
					out<=67;
				end
				if(in == 4) begin
					state<=1965;
					out<=68;
				end
			end
			7745: begin
				if(in == 0) begin
					state<=7756;
					out<=69;
				end
				if(in == 1) begin
					state<=800;
					out<=70;
				end
				if(in == 2) begin
					state<=3867;
					out<=71;
				end
				if(in == 3) begin
					state<=5855;
					out<=72;
				end
				if(in == 4) begin
					state<=1966;
					out<=73;
				end
			end
			7746: begin
				if(in == 0) begin
					state<=7757;
					out<=74;
				end
				if(in == 1) begin
					state<=800;
					out<=75;
				end
				if(in == 2) begin
					state<=3868;
					out<=76;
				end
				if(in == 3) begin
					state<=5856;
					out<=77;
				end
				if(in == 4) begin
					state<=1967;
					out<=78;
				end
			end
			7747: begin
				if(in == 0) begin
					state<=7748;
					out<=79;
				end
				if(in == 1) begin
					state<=800;
					out<=80;
				end
				if(in == 2) begin
					state<=3859;
					out<=81;
				end
				if(in == 3) begin
					state<=5847;
					out<=82;
				end
				if(in == 4) begin
					state<=1958;
					out<=83;
				end
			end
			7748: begin
				if(in == 0) begin
					state<=7759;
					out<=84;
				end
				if(in == 1) begin
					state<=800;
					out<=85;
				end
				if(in == 2) begin
					state<=3870;
					out<=86;
				end
				if(in == 3) begin
					state<=5858;
					out<=87;
				end
				if(in == 4) begin
					state<=1969;
					out<=88;
				end
			end
			7749: begin
				if(in == 0) begin
					state<=7760;
					out<=89;
				end
				if(in == 1) begin
					state<=800;
					out<=90;
				end
				if(in == 2) begin
					state<=3871;
					out<=91;
				end
				if(in == 3) begin
					state<=5859;
					out<=92;
				end
				if(in == 4) begin
					state<=1970;
					out<=93;
				end
			end
			7750: begin
				if(in == 0) begin
					state<=7761;
					out<=94;
				end
				if(in == 1) begin
					state<=800;
					out<=95;
				end
				if(in == 2) begin
					state<=3872;
					out<=96;
				end
				if(in == 3) begin
					state<=5860;
					out<=97;
				end
				if(in == 4) begin
					state<=1971;
					out<=98;
				end
			end
			7751: begin
				if(in == 0) begin
					state<=7762;
					out<=99;
				end
				if(in == 1) begin
					state<=800;
					out<=100;
				end
				if(in == 2) begin
					state<=3873;
					out<=101;
				end
				if(in == 3) begin
					state<=5861;
					out<=102;
				end
				if(in == 4) begin
					state<=1972;
					out<=103;
				end
			end
			7752: begin
				if(in == 0) begin
					state<=7763;
					out<=104;
				end
				if(in == 1) begin
					state<=800;
					out<=105;
				end
				if(in == 2) begin
					state<=3874;
					out<=106;
				end
				if(in == 3) begin
					state<=5862;
					out<=107;
				end
				if(in == 4) begin
					state<=1973;
					out<=108;
				end
			end
			7753: begin
				if(in == 0) begin
					state<=7764;
					out<=109;
				end
				if(in == 1) begin
					state<=800;
					out<=110;
				end
				if(in == 2) begin
					state<=3875;
					out<=111;
				end
				if(in == 3) begin
					state<=5863;
					out<=112;
				end
				if(in == 4) begin
					state<=1974;
					out<=113;
				end
			end
			7754: begin
				if(in == 0) begin
					state<=7765;
					out<=114;
				end
				if(in == 1) begin
					state<=800;
					out<=115;
				end
				if(in == 2) begin
					state<=3876;
					out<=116;
				end
				if(in == 3) begin
					state<=5864;
					out<=117;
				end
				if(in == 4) begin
					state<=1975;
					out<=118;
				end
			end
			7755: begin
				if(in == 0) begin
					state<=7766;
					out<=119;
				end
				if(in == 1) begin
					state<=800;
					out<=120;
				end
				if(in == 2) begin
					state<=3877;
					out<=121;
				end
				if(in == 3) begin
					state<=5865;
					out<=122;
				end
				if(in == 4) begin
					state<=1976;
					out<=123;
				end
			end
			7756: begin
				if(in == 0) begin
					state<=7767;
					out<=124;
				end
				if(in == 1) begin
					state<=800;
					out<=125;
				end
				if(in == 2) begin
					state<=3878;
					out<=126;
				end
				if(in == 3) begin
					state<=5866;
					out<=127;
				end
				if(in == 4) begin
					state<=1977;
					out<=128;
				end
			end
			7757: begin
				if(in == 0) begin
					state<=7758;
					out<=129;
				end
				if(in == 1) begin
					state<=800;
					out<=130;
				end
				if(in == 2) begin
					state<=3869;
					out<=131;
				end
				if(in == 3) begin
					state<=5857;
					out<=132;
				end
				if(in == 4) begin
					state<=1968;
					out<=133;
				end
			end
			7758: begin
				if(in == 0) begin
					state<=7769;
					out<=134;
				end
				if(in == 1) begin
					state<=800;
					out<=135;
				end
				if(in == 2) begin
					state<=3880;
					out<=136;
				end
				if(in == 3) begin
					state<=5868;
					out<=137;
				end
				if(in == 4) begin
					state<=1979;
					out<=138;
				end
			end
			7759: begin
				if(in == 0) begin
					state<=7770;
					out<=139;
				end
				if(in == 1) begin
					state<=800;
					out<=140;
				end
				if(in == 2) begin
					state<=3881;
					out<=141;
				end
				if(in == 3) begin
					state<=5869;
					out<=142;
				end
				if(in == 4) begin
					state<=1980;
					out<=143;
				end
			end
			7760: begin
				if(in == 0) begin
					state<=7771;
					out<=144;
				end
				if(in == 1) begin
					state<=800;
					out<=145;
				end
				if(in == 2) begin
					state<=3882;
					out<=146;
				end
				if(in == 3) begin
					state<=5870;
					out<=147;
				end
				if(in == 4) begin
					state<=1981;
					out<=148;
				end
			end
			7761: begin
				if(in == 0) begin
					state<=7772;
					out<=149;
				end
				if(in == 1) begin
					state<=800;
					out<=150;
				end
				if(in == 2) begin
					state<=3883;
					out<=151;
				end
				if(in == 3) begin
					state<=5871;
					out<=152;
				end
				if(in == 4) begin
					state<=1982;
					out<=153;
				end
			end
			7762: begin
				if(in == 0) begin
					state<=7773;
					out<=154;
				end
				if(in == 1) begin
					state<=800;
					out<=155;
				end
				if(in == 2) begin
					state<=3884;
					out<=156;
				end
				if(in == 3) begin
					state<=5872;
					out<=157;
				end
				if(in == 4) begin
					state<=1983;
					out<=158;
				end
			end
			7763: begin
				if(in == 0) begin
					state<=7774;
					out<=159;
				end
				if(in == 1) begin
					state<=800;
					out<=160;
				end
				if(in == 2) begin
					state<=3885;
					out<=161;
				end
				if(in == 3) begin
					state<=5873;
					out<=162;
				end
				if(in == 4) begin
					state<=1984;
					out<=163;
				end
			end
			7764: begin
				if(in == 0) begin
					state<=7775;
					out<=164;
				end
				if(in == 1) begin
					state<=800;
					out<=165;
				end
				if(in == 2) begin
					state<=3886;
					out<=166;
				end
				if(in == 3) begin
					state<=5874;
					out<=167;
				end
				if(in == 4) begin
					state<=1985;
					out<=168;
				end
			end
			7765: begin
				if(in == 0) begin
					state<=7776;
					out<=169;
				end
				if(in == 1) begin
					state<=800;
					out<=170;
				end
				if(in == 2) begin
					state<=3887;
					out<=171;
				end
				if(in == 3) begin
					state<=5875;
					out<=172;
				end
				if(in == 4) begin
					state<=1986;
					out<=173;
				end
			end
			7766: begin
				if(in == 0) begin
					state<=7777;
					out<=174;
				end
				if(in == 1) begin
					state<=800;
					out<=175;
				end
				if(in == 2) begin
					state<=3888;
					out<=176;
				end
				if(in == 3) begin
					state<=5876;
					out<=177;
				end
				if(in == 4) begin
					state<=1987;
					out<=178;
				end
			end
			7767: begin
				if(in == 0) begin
					state<=7768;
					out<=179;
				end
				if(in == 1) begin
					state<=800;
					out<=180;
				end
				if(in == 2) begin
					state<=3879;
					out<=181;
				end
				if(in == 3) begin
					state<=5867;
					out<=182;
				end
				if(in == 4) begin
					state<=1978;
					out<=183;
				end
			end
			7768: begin
				if(in == 0) begin
					state<=7779;
					out<=184;
				end
				if(in == 1) begin
					state<=800;
					out<=185;
				end
				if(in == 2) begin
					state<=3890;
					out<=186;
				end
				if(in == 3) begin
					state<=5878;
					out<=187;
				end
				if(in == 4) begin
					state<=1989;
					out<=188;
				end
			end
			7769: begin
				if(in == 0) begin
					state<=7780;
					out<=189;
				end
				if(in == 1) begin
					state<=800;
					out<=190;
				end
				if(in == 2) begin
					state<=3891;
					out<=191;
				end
				if(in == 3) begin
					state<=5879;
					out<=192;
				end
				if(in == 4) begin
					state<=1990;
					out<=193;
				end
			end
			7770: begin
				if(in == 0) begin
					state<=7781;
					out<=194;
				end
				if(in == 1) begin
					state<=800;
					out<=195;
				end
				if(in == 2) begin
					state<=3892;
					out<=196;
				end
				if(in == 3) begin
					state<=5880;
					out<=197;
				end
				if(in == 4) begin
					state<=1991;
					out<=198;
				end
			end
			7771: begin
				if(in == 0) begin
					state<=7782;
					out<=199;
				end
				if(in == 1) begin
					state<=800;
					out<=200;
				end
				if(in == 2) begin
					state<=3893;
					out<=201;
				end
				if(in == 3) begin
					state<=5881;
					out<=202;
				end
				if(in == 4) begin
					state<=1992;
					out<=203;
				end
			end
			7772: begin
				if(in == 0) begin
					state<=7783;
					out<=204;
				end
				if(in == 1) begin
					state<=800;
					out<=205;
				end
				if(in == 2) begin
					state<=3894;
					out<=206;
				end
				if(in == 3) begin
					state<=5882;
					out<=207;
				end
				if(in == 4) begin
					state<=1993;
					out<=208;
				end
			end
			7773: begin
				if(in == 0) begin
					state<=7784;
					out<=209;
				end
				if(in == 1) begin
					state<=800;
					out<=210;
				end
				if(in == 2) begin
					state<=3895;
					out<=211;
				end
				if(in == 3) begin
					state<=5883;
					out<=212;
				end
				if(in == 4) begin
					state<=1994;
					out<=213;
				end
			end
			7774: begin
				if(in == 0) begin
					state<=7785;
					out<=214;
				end
				if(in == 1) begin
					state<=800;
					out<=215;
				end
				if(in == 2) begin
					state<=3896;
					out<=216;
				end
				if(in == 3) begin
					state<=5884;
					out<=217;
				end
				if(in == 4) begin
					state<=1995;
					out<=218;
				end
			end
			7775: begin
				if(in == 0) begin
					state<=7786;
					out<=219;
				end
				if(in == 1) begin
					state<=800;
					out<=220;
				end
				if(in == 2) begin
					state<=3897;
					out<=221;
				end
				if(in == 3) begin
					state<=5885;
					out<=222;
				end
				if(in == 4) begin
					state<=1996;
					out<=223;
				end
			end
			7776: begin
				if(in == 0) begin
					state<=7787;
					out<=224;
				end
				if(in == 1) begin
					state<=800;
					out<=225;
				end
				if(in == 2) begin
					state<=3898;
					out<=226;
				end
				if(in == 3) begin
					state<=5886;
					out<=227;
				end
				if(in == 4) begin
					state<=1997;
					out<=228;
				end
			end
			7777: begin
				if(in == 0) begin
					state<=7778;
					out<=229;
				end
				if(in == 1) begin
					state<=800;
					out<=230;
				end
				if(in == 2) begin
					state<=3889;
					out<=231;
				end
				if(in == 3) begin
					state<=5877;
					out<=232;
				end
				if(in == 4) begin
					state<=1988;
					out<=233;
				end
			end
			7778: begin
				if(in == 0) begin
					state<=6165;
					out<=234;
				end
				if(in == 1) begin
					state<=800;
					out<=235;
				end
				if(in == 2) begin
					state<=2276;
					out<=236;
				end
				if(in == 3) begin
					state<=4798;
					out<=237;
				end
				if(in == 4) begin
					state<=900;
					out<=238;
				end
			end
			7779: begin
				if(in == 0) begin
					state<=6166;
					out<=239;
				end
				if(in == 1) begin
					state<=800;
					out<=240;
				end
				if(in == 2) begin
					state<=2277;
					out<=241;
				end
				if(in == 3) begin
					state<=4799;
					out<=242;
				end
				if(in == 4) begin
					state<=901;
					out<=243;
				end
			end
			7780: begin
				if(in == 0) begin
					state<=6167;
					out<=244;
				end
				if(in == 1) begin
					state<=800;
					out<=245;
				end
				if(in == 2) begin
					state<=2278;
					out<=246;
				end
				if(in == 3) begin
					state<=4800;
					out<=247;
				end
				if(in == 4) begin
					state<=902;
					out<=248;
				end
			end
			7781: begin
				if(in == 0) begin
					state<=6168;
					out<=249;
				end
				if(in == 1) begin
					state<=800;
					out<=250;
				end
				if(in == 2) begin
					state<=2279;
					out<=251;
				end
				if(in == 3) begin
					state<=4801;
					out<=252;
				end
				if(in == 4) begin
					state<=903;
					out<=253;
				end
			end
			7782: begin
				if(in == 0) begin
					state<=6169;
					out<=254;
				end
				if(in == 1) begin
					state<=800;
					out<=255;
				end
				if(in == 2) begin
					state<=2280;
					out<=0;
				end
				if(in == 3) begin
					state<=4802;
					out<=1;
				end
				if(in == 4) begin
					state<=904;
					out<=2;
				end
			end
			7783: begin
				if(in == 0) begin
					state<=6170;
					out<=3;
				end
				if(in == 1) begin
					state<=800;
					out<=4;
				end
				if(in == 2) begin
					state<=2281;
					out<=5;
				end
				if(in == 3) begin
					state<=4803;
					out<=6;
				end
				if(in == 4) begin
					state<=905;
					out<=7;
				end
			end
			7784: begin
				if(in == 0) begin
					state<=6171;
					out<=8;
				end
				if(in == 1) begin
					state<=800;
					out<=9;
				end
				if(in == 2) begin
					state<=2282;
					out<=10;
				end
				if(in == 3) begin
					state<=4804;
					out<=11;
				end
				if(in == 4) begin
					state<=906;
					out<=12;
				end
			end
			7785: begin
				if(in == 0) begin
					state<=6172;
					out<=13;
				end
				if(in == 1) begin
					state<=800;
					out<=14;
				end
				if(in == 2) begin
					state<=2283;
					out<=15;
				end
				if(in == 3) begin
					state<=4805;
					out<=16;
				end
				if(in == 4) begin
					state<=907;
					out<=17;
				end
			end
			7786: begin
				if(in == 0) begin
					state<=6173;
					out<=18;
				end
				if(in == 1) begin
					state<=800;
					out<=19;
				end
				if(in == 2) begin
					state<=2284;
					out<=20;
				end
				if(in == 3) begin
					state<=4806;
					out<=21;
				end
				if(in == 4) begin
					state<=908;
					out<=22;
				end
			end
			7787: begin
				if(in == 0) begin
					state<=6164;
					out<=23;
				end
				if(in == 1) begin
					state<=800;
					out<=24;
				end
				if(in == 2) begin
					state<=2275;
					out<=25;
				end
				if(in == 3) begin
					state<=5887;
					out<=26;
				end
				if(in == 4) begin
					state<=1998;
					out<=27;
				end
			end
		endcase
	end
endmodule